-- @file rom_font.vhd
-- @brief ROM containing character font
-- @author Justin Davis
--
-- $Revision: -
-- $Date: 06/22/2023
-- $LastEditedBy: Justin Davis
--
-- Developed by 2023 Southwest Research Institute
-------------------------------------------------------------------------------
-- Font data taken from: https://github.com/robhagemans/hoard-of-bitfonts/blob/master/atari/8-bit/atascii.yaff

library ieee;           use ieee.std_logic_1164.all;
                        use ieee.numeric_std.all;

library work;           use work.tools_pkg.all;
                        use work.sys_description_pkg.all;

entity rom_font is
    port ( addrIn   : in    slv(10 downto 0) ;
           dataOut  :   out slv(7 downto 0));
end entity rom_font;

architecture rtl of rom_font is
   
    type rom_type is array (0 to (2**addrIn'length)-1) of std_logic_vector(dataOut'range);

	-- ROM definition
    signal rom : rom_type := ( 

-- # [?] BLACK HEART SUIT
-- u+2665:
-- 0x00:
    "00000000",
    "00110110",
    "01111111",
    "01111111",
    "00111110",
    "00011100",
    "00001000",
    "00000000",


-- # [?] BOX DRAWINGS LIGHT VERTICAL AND RIGHT
-- u+251c:
-- 0x01:
    "00011000",
    "00011000",
    "00011000",
    "00011111",
    "00011111",
    "00011000",
    "00011000",
    "00011000",


-- # [?] RIGHT VERTICAL BOX LINE
-- u+23b9:
-- 0x02:
    "00000011",
    "00000011",
    "00000011",
    "00000011",
    "00000011",
    "00000011",
    "00000011",
    "00000011",


-- # [?] BOX DRAWINGS LIGHT UP AND LEFT
-- u+2518:
-- 0x03:
    "00011000",
    "00011000",
    "00011000",
    "11111000",
    "11111000",
    "00000000",
    "00000000",
    "00000000",


-- # [?] BOX DRAWINGS LIGHT VERTICAL AND LEFT
-- u+2524:
-- 0x04:
    "00011000",
    "00011000",
    "00011000",
    "11111000",
    "11111000",
    "00011000",
    "00011000",
    "00011000",


-- # [?] BOX DRAWINGS LIGHT DOWN AND LEFT
-- u+2510:
-- 0x05:
    "00000000",
    "00000000",
    "00000000",
    "11111000",
    "11111000",
    "00011000",
    "00011000",
    "00011000",


-- # [?] BOX DRAWINGS LIGHT DIAGONAL UPPER RIGHT TO LOWER LEFT
-- u+2571:
-- 0x06:
    "00000011",
    "00000111",
    "00001110",
    "00011100",
    "00111000",
    "01110000",
    "11100000",
    "11000000",


-- # [?] BOX DRAWINGS LIGHT DIAGONAL UPPER LEFT TO LOWER RIGHT
-- u+2572:
-- 0x07:
    "11000000",
    "11100000",
    "01110000",
    "00111000",
    "00011100",
    "00001110",
    "00000111",
    "00000011",


-- # [?] BLACK LOWER RIGHT TRIANGLE
-- u+25e2:
-- 0x08:
    "00000001",
    "00000011",
    "00000111",
    "00001111",
    "00011111",
    "00111111",
    "01111111",
    "11111111",


-- # [?] QUADRANT LOWER RIGHT
-- u+2597:
-- 0x09:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00001111",
    "00001111",
    "00001111",
    "00001111",


-- # [?] BLACK LOWER LEFT TRIANGLE
-- u+25e3:
-- 0x0a:
    "10000000",
    "11000000",
    "11100000",
    "11110000",
    "11111000",
    "11111100",
    "11111110",
    "11111111",


-- # [?] QUADRANT UPPER RIGHT
-- u+259d:
-- 0x0b:
    "00001111",
    "00001111",
    "00001111",
    "00001111",
    "00000000",
    "00000000",
    "00000000",
    "00000000",


-- # [?] QUADRANT UPPER LEFT
-- u+2598:
-- 0x0c:
    "11110000",
    "11110000",
    "11110000",
    "11110000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",


-- # [?] HORIZONTAL SCAN LINE-1",
-- u+23ba:
-- 0x0d:
    "11111111",
    "11111111",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",


-- # [?] HORIZONTAL SCAN LINE-9
-- u+23bd:
-- 0x0e:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111111",
    "11111111",


-- # [?] QUADRANT LOWER LEFT
-- u+2596:
-- 0x0f:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11110000",
    "11110000",
    "11110000",
    "11110000",


-- # [?] BLACK CLUB SUIT
-- u+2663:
-- 0x10:
    "00000000",
    "00011100",
    "00011100",
    "01110111",
    "01110111",
    "00001000",
    "00011100",
    "00000000",


-- # [?] BOX DRAWINGS LIGHT DOWN AND RIGHT
-- u+250c:
-- 0x11:
    "00000000",
    "00000000",
    "00000000",
    "00011111",
    "00011111",
    "00011000",
    "00011000",
    "00011000",


-- # [?] BOX DRAWINGS LIGHT HORIZONTAL
-- u+2500:
-- 0x12:
    "00000000",
    "00000000",
    "00000000",
    "11111111",
    "11111111",
    "00000000",
    "00000000",
    "00000000",


-- # [?] BOX DRAWINGS LIGHT VERTICAL AND HORIZONTAL
-- u+253c:
-- 0x13:
    "00011000",
    "00011000",
    "00011000",
    "11111111",
    "11111111",
    "00011000",
    "00011000",
    "00011000",


-- # [�] BULLET
-- u+2022:
-- 0x14:
    "00000000",
    "00000000",
    "00111100",
    "01111110",
    "01111110",
    "01111110",
    "00111100",
    "00000000",


-- # [?] LOWER HALF BLOCK
-- u+2584:
-- 0x15:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111111",
    "11111111",
    "11111111",
    "11111111",


-- # [?] LEFT VERTICAL BOX LINE
-- u+23b8:
-- 0x16:
    "11000000",
    "11000000",
    "11000000",
    "11000000",
    "11000000",
    "11000000",
    "11000000",
    "11000000",


-- # [?] BOX DRAWINGS LIGHT DOWN AND HORIZONTAL
-- u+252c:
-- 0x17:
    "00000000",
    "00000000",
    "00000000",
    "11111111",
    "11111111",
    "00011000",
    "00011000",
    "00011000",


-- # [?] BOX DRAWINGS LIGHT UP AND HORIZONTAL
-- u+2534:
-- 0x18:
    "00011000",
    "00011000",
    "00011000",
    "11111111",
    "11111111",
    "00000000",
    "00000000",
    "00000000",


-- # [?] LEFT HALF BLOCK
-- u+258c:
-- 0x19:
    "11110000",
    "11110000",
    "11110000",
    "11110000",
    "11110000",
    "11110000",
    "11110000",
    "11110000",


-- # [?] BOX DRAWINGS LIGHT UP AND RIGHT
-- u+2514:
-- 0x1a:
    "00011000",
    "00011000",
    "00011000",
    "00011111",
    "00011111",
    "00000000",
    "00000000",
    "00000000",

-- 0x1b:
    "01111000",
    "01100000",
    "01111000",
    "01100000",
    "01111110",
    "00011000",
    "00011110",
    "00000000",

-- 0x1c:
    "00000000",
    "00011000",
    "00111100",
    "01111110",
    "00011000",
    "00011000",
    "00011000",
    "00000000",

-- 0x1d:
    "00000000",
    "00011000",
    "00011000",
    "00011000",
    "01111110",
    "00111100",
    "00011000",
    "00000000",

-- 0x1e:
    "00000000",
    "00011000",
    "00110000",
    "01111110",
    "00110000",
    "00011000",
    "00000000",
    "00000000",

-- 0x1f:
    "00000000",
    "00011000",
    "00001100",
    "01111110",
    "00001100",
    "00011000",
    "00000000",
    "00000000",


-- # [ ] SPACE
-- u+0020:
-- 0x20:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",


-- # [!] EXCLAMATION MARK
-- u+0021:
-- 0x21:
    "00000000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00000000",
    "00011000",
    "00000000",


-- # ["] QUOTATION MARK
-- u+0022:
-- 0x22:
    "00000000",
    "01100110",
    "01100110",
    "01100110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",


-- # [-- #] NUMBER SIGN
-- u+0023:
-- 0x23:
    "00000000",
    "01100110",
    "11111111",
    "01100110",
    "01100110",
    "11111111",
    "01100110",
    "00000000",


-- # [$] DOLLAR SIGN
-- u+0024:
-- 0x24:
    "00011000",
    "00111110",
    "01100000",
    "00111100",
    "00000110",
    "01111100",
    "00011000",
    "00000000",


-- # [%] PERCENT SIGN
-- u+0025:
-- 0x25:
    "00000000",
    "01100110",
    "01101100",
    "00011000",
    "00110000",
    "01100110",
    "01000110",
    "00000000",


-- # [&] AMPERSAND
-- u+0026:
-- 0x26:
    "00011100",
    "00110110",
    "00011100",
    "00111000",
    "01101111",
    "01100110",
    "00111011",
    "00000000",


-- # ['] APOSTROPHE
-- u+0027:
-- 0x27:
    "00000000",
    "00011000",
    "00011000",
    "00011000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",


-- # [(] LEFT PARENTHESIS
-- u+0028:
-- 0x28:
    "00000000",
    "00001110",
    "00011100",
    "00011000",
    "00011000",
    "00011100",
    "00001110",
    "00000000",


-- # [)] RIGHT PARENTHESIS
-- u+0029:
-- 0x29:
    "00000000",
    "01110000",
    "00111000",
    "00011000",
    "00011000",
    "00111000",
    "01110000",
    "00000000",


-- # [*] ASTERISK
-- u+002a:
-- 0x2a:
    "00000000",
    "01100110",
    "00111100",
    "11111111",
    "00111100",
    "01100110",
    "00000000",
    "00000000",


-- # [+] PLUS SIGN
-- u+002b:
-- 0x2b:
    "00000000",
    "00011000",
    "00011000",
    "01111110",
    "00011000",
    "00011000",
    "00000000",
    "00000000",


-- # [,] COMMA
-- u+002c:
-- 0x2c:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011000",
    "00011000",
    "00110000",


-- # [-] HYPHEN-MINUS
-- u+002d:
-- 0x2d:
    "00000000",
    "00000000",
    "00000000",
    "01111110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",


-- # [0] FULL STOP
-- u+002e:
-- 0x2e:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011000",
    "00011000",
    "00000000",


-- # [/] SOLIDUS
-- u+002f:
-- 0x2f:
    "00000000",
    "00000110",
    "00001100",
    "00011000",
    "00110000",
    "01100000",
    "01000000",
    "00000000",


-- # [0] DIGIT ZERO
-- u+0030:
-- 0x30:
    "00000000",
    "00111100",
    "01100110",
    "01101110",
    "01110110",
    "01100110",
    "00111100",
    "00000000",


-- # [1] DIGIT ONE
-- u+0031:
-- 0x31:
    "00000000",
    "00011000",
    "00111000",
    "00011000",
    "00011000",
    "00011000",
    "01111110",
    "00000000",


-- # [2] DIGIT TWO
-- u+0032:
-- 0x32:
    "00000000",
    "00111100",
    "01100110",
    "00001100",
    "00011000",
    "00110000",
    "01111110",
    "00000000",


-- # [3] DIGIT THREE
-- u+0033:
-- 0x33:
    "00000000",
    "01111110",
    "00001100",
    "00011000",
    "00001100",
    "01100110",
    "00111100",
    "00000000",


-- # [4] DIGIT FOUR
-- u+0034:
-- 0x34:
    "00000000",
    "00001100",
    "00011100",
    "00111100",
    "01101100",
    "01111110",
    "00001100",
    "00000000",


-- # [5] DIGIT FIVE
-- u+0035:
-- 0x35:
    "00000000",
    "01111110",
    "01100000",
    "01111100",
    "00000110",
    "01100110",
    "00111100",
    "00000000",


-- # [6] DIGIT SIX
-- u+0036:
-- 0x36:
    "00000000",
    "00111100",
    "01100000",
    "01111100",
    "01100110",
    "01100110",
    "00111100",
    "00000000",


-- # [7] DIGIT SEVEN
-- u+0037:
-- 0x37:
    "00000000",
    "01111110",
    "00000110",
    "00001100",
    "00011000",
    "00110000",
    "00110000",
    "00000000",


-- # [8] DIGIT EIGHT
-- u+0038:
-- 0x38:
    "00000000",
    "00111100",
    "01100110",
    "00111100",
    "01100110",
    "01100110",
    "00111100",
    "00000000",


-- # [9] DIGIT NINE
-- u+0039:
-- 0x39:
    "00000000",
    "00111100",
    "01100110",
    "00111110",
    "00000110",
    "00001100",
    "00111000",
    "00000000",


-- # [:] COLON
-- u+003a:
-- 0x3a:
    "00000000",
    "00000000",
    "00011000",
    "00011000",
    "00000000",
    "00011000",
    "00011000",
    "00000000",


-- # [;] SEMICOLON
-- u+003b:
-- 0x3b:
    "00000000",
    "00000000",
    "00011000",
    "00011000",
    "00000000",
    "00011000",
    "00011000",
    "00110000",


-- # [<] LESS-THAN SIGN
-- u+003c:
-- 0x3c:
    "00000110",
    "00001100",
    "00011000",
    "00110000",
    "00011000",
    "00001100",
    "00000110",
    "00000000",


-- # [=] EQUALS SIGN
-- u+003d:
-- 0x3d:
    "00000000",
    "00000000",
    "01111110",
    "00000000",
    "00000000",
    "01111110",
    "00000000",
    "00000000",


-- # [>] GREATER-THAN SIGN
-- u+003e:
-- 0x3e:
    "01100000",
    "00110000",
    "00011000",
    "00001100",
    "00011000",
    "00110000",
    "01100000",
    "00000000",


-- # [?] QUESTION MARK
-- u+003f:
-- 0x3f:
    "00000000",
    "00111100",
    "01100110",
    "00001100",
    "00011000",
    "00000000",
    "00011000",
    "00000000",


-- # [1] COMMERCIAL AT
-- u+0040:
-- 0x40:
    "00000000",
    "00111100",
    "01100110",
    "01101110",
    "01101110",
    "01100000",
    "00111110",
    "00000000",


-- # [A] LATIN CAPITAL LETTER A
-- u+0041:
-- 0x41:
    "00000000",
    "00011000",
    "00111100",
    "01100110",
    "01100110",
    "01111110",
    "01100110",
    "00000000",


-- # [B] LATIN CAPITAL LETTER B
-- u+0042:
-- 0x42:
    "00000000",
    "01111100",
    "01100110",
    "01111100",
    "01100110",
    "01100110",
    "01111100",
    "00000000",


-- # [C] LATIN CAPITAL LETTER C
-- u+0043:
-- 0x43:
    "00000000",
    "00111100",
    "01100110",
    "01100000",
    "01100000",
    "01100110",
    "00111100",
    "00000000",


-- # [D] LATIN CAPITAL LETTER D
-- u+0044:
-- 0x44:
    "00000000",
    "01111000",
    "01101100",
    "01100110",
    "01100110",
    "01101100",
    "01111000",
    "00000000",


-- # [E] LATIN CAPITAL LETTER E
-- u+0045:
-- 0x45:
    "00000000",
    "01111110",
    "01100000",
    "01111100",
    "01100000",
    "01100000",
    "01111110",
    "00000000",


-- # [F] LATIN CAPITAL LETTER F
-- u+0046:
-- 0x46:
    "00000000",
    "01111110",
    "01100000",
    "01111100",
    "01100000",
    "01100000",
    "01100000",
    "00000000",


-- # [G] LATIN CAPITAL LETTER G
-- u+0047:
-- 0x47:
    "00000000",
    "00111110",
    "01100000",
    "01100000",
    "01101110",
    "01100110",
    "00111110",
    "00000000",


-- # [H] LATIN CAPITAL LETTER H
-- u+0048:
-- 0x48:
    "00000000",
    "01100110",
    "01100110",
    "01111110",
    "01100110",
    "01100110",
    "01100110",
    "00000000",


-- # [I] LATIN CAPITAL LETTER I
-- u+0049:
-- 0x49:
    "00000000",
    "01111110",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "01111110",
    "00000000",


-- # [J] LATIN CAPITAL LETTER J
-- u+004a:
-- 0x4a:
    "00000000",
    "00000110",
    "00000110",
    "00000110",
    "00000110",
    "01100110",
    "00111100",
    "00000000",


-- # [K] LATIN CAPITAL LETTER K
-- u+004b:
-- 0x4b:
    "00000000",
    "01100110",
    "01101100",
    "01111000",
    "01111000",
    "01101100",
    "01100110",
    "00000000",


-- # [L] LATIN CAPITAL LETTER L
-- u+004c:
-- 0x4c:
    "00000000",
    "01100000",
    "01100000",
    "01100000",
    "01100000",
    "01100000",
    "01111110",
    "00000000",


-- # [M] LATIN CAPITAL LETTER M
-- u+004d:
-- 0x4d:
    "00000000",
    "01100011",
    "01110111",
    "01111111",
    "01101011",
    "01100011",
    "01100011",
    "00000000",


-- # [N] LATIN CAPITAL LETTER N
-- u+004e:
-- 0x4e:
    "00000000",
    "01100110",
    "01110110",
    "01111110",
    "01111110",
    "01101110",
    "01100110",
    "00000000",


-- # [O] LATIN CAPITAL LETTER O
-- u+004f:
-- 0x4f:
    "00000000",
    "00111100",
    "01100110",
    "01100110",
    "01100110",
    "01100110",
    "00111100",
    "00000000",


-- # [P] LATIN CAPITAL LETTER P
-- u+0050:
-- 0x50:
    "00000000",
    "01111100",
    "01100110",
    "01100110",
    "01111100",
    "01100000",
    "01100000",
    "00000000",


-- # [Q] LATIN CAPITAL LETTER Q
-- u+0051:
-- 0x51:
    "00000000",
    "00111100",
    "01100110",
    "01100110",
    "01100110",
    "01101100",
    "00110110",
    "00000000",


-- # [R] LATIN CAPITAL LETTER R
-- u+0052:
-- 0x52:
    "00000000",
    "01111100",
    "01100110",
    "01100110",
    "01111100",
    "01101100",
    "01100110",
    "00000000",


-- # [S] LATIN CAPITAL LETTER S
-- u+0053:
-- 0x53:
    "00000000",
    "00111100",
    "01100000",
    "00111100",
    "00000110",
    "00000110",
    "00111100",
    "00000000",


-- # [T] LATIN CAPITAL LETTER T
-- u+0054:
-- 0x54:
    "00000000",
    "01111110",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00000000",


-- # [U] LATIN CAPITAL LETTER U
-- u+0055:
-- 0x55:
    "00000000",
    "01100110",
    "01100110",
    "01100110",
    "01100110",
    "01100110",
    "01111110",
    "00000000",


-- # [V] LATIN CAPITAL LETTER V
-- u+0056:
-- 0x56:
    "00000000",
    "01100110",
    "01100110",
    "01100110",
    "01100110",
    "00111100",
    "00011000",
    "00000000",


-- # [W] LATIN CAPITAL LETTER W
-- u+0057:
-- 0x57:
    "00000000",
    "01100011",
    "01100011",
    "01101011",
    "01111111",
    "01110111",
    "01100011",
    "00000000",


-- # [X] LATIN CAPITAL LETTER X
-- u+0058:
-- 0x58:
    "00000000",
    "01100110",
    "01100110",
    "00111100",
    "00111100",
    "01100110",
    "01100110",
    "00000000",


-- # [Y] LATIN CAPITAL LETTER Y
-- u+0059:
-- 0x59:
    "00000000",
    "01100110",
    "01100110",
    "00111100",
    "00011000",
    "00011000",
    "00011000",
    "00000000",


-- # [Z] LATIN CAPITAL LETTER Z
-- u+005a:
-- 0x5a:
    "00000000",
    "01111110",
    "00001100",
    "00011000",
    "00110000",
    "01100000",
    "01111110",
    "00000000",


-- # [[] LEFT SQUARE BRACKET
-- u+005b:
-- 0x5b:
    "00000000",
    "00011110",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011110",
    "00000000",


-- # [\] REVERSE SOLIDUS
-- u+005c:
-- 0x5c:
    "00000000",
    "01000000",
    "01100000",
    "00110000",
    "00011000",
    "00001100",
    "00000110",
    "00000000",


-- # []] RIGHT SQUARE BRACKET
-- u+005d:
-- 0x5d:
    "00000000",
    "01111000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "01111000",
    "00000000",


-- # [^] CIRCUMFLEX ACCENT
-- u+005e:
-- 0x5e:
    "00000000",
    "00001000",
    "00011100",
    "00110110",
    "01100011",
    "00000000",
    "00000000",
    "00000000",


-- # [_] LOW LINE
-- u+005f:
-- 0x5f:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111111",
    "00000000",


-- # [?] BLACK DIAMOND SUIT
-- u+2666:
-- 0x60:
    "00000000",
    "00011000",
    "00111100",
    "01111110",
    "01111110",
    "00111100",
    "00011000",
    "00000000",


-- # [a] LATIN SMALL LETTER A
-- u+0061:
-- 0x61:
    "00000000",
    "00000000",
    "00111100",
    "00000110",
    "00111110",
    "01100110",
    "00111110",
    "00000000",


-- # [b] LATIN SMALL LETTER B
-- u+0062:
-- 0x62:
    "00000000",
    "01100000",
    "01100000",
    "01111100",
    "01100110",
    "01100110",
    "01111100",
    "00000000",


-- # [c] LATIN SMALL LETTER C
-- u+0063:
-- 0x63:
    "00000000",
    "00000000",
    "00111100",
    "01100000",
    "01100000",
    "01100000",
    "00111100",
    "00000000",


-- # [d] LATIN SMALL LETTER D
-- u+0064:
-- 0x64:
    "00000000",
    "00000110",
    "00000110",
    "00111110",
    "01100110",
    "01100110",
    "00111110",
    "00000000",


-- # [e] LATIN SMALL LETTER E
-- u+0065:
-- 0x65:
    "00000000",
    "00000000",
    "00111100",
    "01100110",
    "01111110",
    "01100000",
    "00111100",
    "00000000",


-- # [f] LATIN SMALL LETTER F
-- u+0066:
-- 0x66:
    "00000000",
    "00001110",
    "00011000",
    "00111110",
    "00011000",
    "00011000",
    "00011000",
    "00000000",


-- # [g] LATIN SMALL LETTER G
-- u+0067:
-- 0x67:
    "00000000",
    "00000000",
    "00111110",
    "01100110",
    "01100110",
    "00111110",
    "00000110",
    "01111100",


-- # [h] LATIN SMALL LETTER H
-- u+0068:
-- 0x68:
    "00000000",
    "01100000",
    "01100000",
    "01111100",
    "01100110",
    "01100110",
    "01100110",
    "00000000",


-- # [i] LATIN SMALL LETTER I
-- u+0069:
-- 0x69:
    "00000000",
    "00011000",
    "00000000",
    "00111000",
    "00011000",
    "00011000",
    "00111100",
    "00000000",


-- # [j] LATIN SMALL LETTER J
-- u+006a:
-- 0x6a:
    "00000000",
    "00000110",
    "00000000",
    "00000110",
    "00000110",
    "00000110",
    "00000110",
    "00111100",


-- # [k] LATIN SMALL LETTER K
-- u+006b:
-- 0x6b:
    "00000000",
    "01100000",
    "01100000",
    "01101100",
    "01111000",
    "01101100",
    "01100110",
    "00000000",


-- # [l] LATIN SMALL LETTER L
-- u+006c:
-- 0x6c:
    "00000000",
    "00111000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00111100",
    "00000000",


-- # [m] LATIN SMALL LETTER M
-- u+006d:
-- 0x6d:
    "00000000",
    "00000000",
    "01100110",
    "01111111",
    "01111111",
    "01101011",
    "01100011",
    "00000000",


-- # [n] LATIN SMALL LETTER N
-- u+006e:
-- 0x6e:
    "00000000",
    "00000000",
    "01111100",
    "01100110",
    "01100110",
    "01100110",
    "01100110",
    "00000000",


-- # [o] LATIN SMALL LETTER O
-- u+006f:
-- 0x6f:
    "00000000",
    "00000000",
    "00111100",
    "01100110",
    "01100110",
    "01100110",
    "00111100",
    "00000000",


-- # [p] LATIN SMALL LETTER P
-- u+0070:
-- 0x70:
    "00000000",
    "00000000",
    "01111100",
    "01100110",
    "01100110",
    "01111100",
    "01100000",
    "01100000",


-- # [q] LATIN SMALL LETTER Q
-- u+0071:
-- 0x71:
    "00000000",
    "00000000",
    "00111110",
    "01100110",
    "01100110",
    "00111110",
    "00000110",
    "00000110",


-- # [r] LATIN SMALL LETTER R
-- u+0072:
-- 0x72:
    "00000000",
    "00000000",
    "01111100",
    "01100110",
    "01100000",
    "01100000",
    "01100000",
    "00000000",


-- # [s] LATIN SMALL LETTER S
-- u+0073:
-- 0x73:
    "00000000",
    "00000000",
    "00111110",
    "01100000",
    "00111100",
    "00000110",
    "01111100",
    "00000000",


-- # [t] LATIN SMALL LETTER T
-- u+0074:
-- 0x74:
    "00000000",
    "00011000",
    "01111110",
    "00011000",
    "00011000",
    "00011000",
    "00001110",
    "00000000",


-- # [u] LATIN SMALL LETTER U
-- u+0075:
-- 0x75:
    "00000000",
    "00000000",
    "01100110",
    "01100110",
    "01100110",
    "01100110",
    "00111110",
    "00000000",


-- # [v] LATIN SMALL LETTER V
-- u+0076:
-- 0x76:
    "00000000",
    "00000000",
    "01100110",
    "01100110",
    "01100110",
    "00111100",
    "00011000",
    "00000000",


-- # [w] LATIN SMALL LETTER W
-- u+0077:
-- 0x77:
    "00000000",
    "00000000",
    "01100011",
    "01101011",
    "01111111",
    "00111110",
    "00110110",
    "00000000",


-- # [x] LATIN SMALL LETTER X
-- u+0078:
-- 0x78:
    "00000000",
    "00000000",
    "01100110",
    "00111100",
    "00011000",
    "00111100",
    "01100110",
    "00000000",


-- # [y] LATIN SMALL LETTER Y
-- u+0079:
-- 0x79:
    "00000000",
    "00000000",
    "01100110",
    "01100110",
    "01100110",
    "00111110",
    "00001100",
    "01111000",


-- # [z] LATIN SMALL LETTER Z
-- u+007a:
-- 0x7a:
    "00000000",
    "00000000",
    "01111110",
    "00001100",
    "00011000",
    "00110000",
    "01111110",
    "00000000",


-- # [?] BLACK SPADE SUIT
-- u+2660:
-- 0x7b:
    "00000000",
    "00011000",
    "00111100",
    "01111110",
    "01111110",
    "00011000",
    "00111100",
    "00000000",


-- # [|] VERTICAL LINE
-- u+007c:
-- 0x7c:
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",
    "00011000",

-- 0x7d:
    "00000000",
    "01111110",
    "01111000",
    "01111100",
    "01101110",
    "01100110",
    "00000110",
    "00000000",

-- 0x7e:
    "00001000",
    "00011000",
    "00111000",
    "01111000",
    "00111000",
    "00011000",
    "00001000",
    "00000000",

-- 0x7f:
    "00010000",
    "00011000",
    "00011100",
    "00011110",
    "00011100",
    "00011000",
    "00010000",
    "00000000",


-- # [?] BLACK HEART SUIT
-- u+2665:
-- 0x80:
    "11111111",
    "11001001",
    "10000000",
    "10000000",
    "11000001",
    "11100011",
    "11110111",
    "11111111",


-- # [?] BOX DRAWINGS LIGHT VERTICAL AND RIGHT
-- u+251c:
-- 0x81:
    "11100111",
    "11100111",
    "11100111",
    "11100000",
    "11100000",
    "11100111",
    "11100111",
    "11100111",


-- # [?] RIGHT VERTICAL BOX LINE
-- u+23b9:
-- 0x82:
    "11111100",
    "11111100",
    "11111100",
    "11111100",
    "11111100",
    "11111100",
    "11111100",
    "11111100",


-- # [?] BOX DRAWINGS LIGHT UP AND LEFT
-- u+2518:
-- 0x83:
    "11100111",
    "11100111",
    "11100111",
    "00000111",
    "00000111",
    "11111111",
    "11111111",
    "11111111",


-- # [?] BOX DRAWINGS LIGHT VERTICAL AND LEFT
-- u+2524:
-- 0x84:
    "11100111",
    "11100111",
    "11100111",
    "00000111",
    "00000111",
    "11100111",
    "11100111",
    "11100111",


-- # [?] BOX DRAWINGS LIGHT DOWN AND LEFT
-- u+2510:
-- 0x85:
    "11111111",
    "11111111",
    "11111111",
    "00000111",
    "00000111",
    "11100111",
    "11100111",
    "11100111",


-- # [?] BOX DRAWINGS LIGHT DIAGONAL UPPER RIGHT TO LOWER LEFT
-- u+2571:
-- 0x86:
    "11111100",
    "11111000",
    "11110001",
    "11100011",
    "11000111",
    "10001111",
    "00011111",
    "00111111",


-- # [?] BOX DRAWINGS LIGHT DIAGONAL UPPER LEFT TO LOWER RIGHT
-- u+2572:
-- 0x87:
    "00111111",
    "00011111",
    "10001111",
    "11000111",
    "11100011",
    "11110001",
    "11111000",
    "11111100",


-- # [?] BLACK UPPER LEFT TRIANGLE
-- u+25e4:
-- 0x88:
    "11111110",
    "11111100",
    "11111000",
    "11110000",
    "11100000",
    "11000000",
    "10000000",
    "00000000",


-- # [?] QUADRANT UPPER LEFT AND UPPER RIGHT AND LOWER LEFT
-- u+259b:
-- 0x89:
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11110000",
    "11110000",
    "11110000",
    "11110000",


-- # [?] BLACK UPPER RIGHT TRIANGLE
-- u+25e5:
-- 0x8a:
    "01111111",
    "00111111",
    "00011111",
    "00001111",
    "00000111",
    "00000011",
    "00000001",
    "00000000",


-- # [?] QUADRANT UPPER LEFT AND LOWER LEFT AND LOWER RIGHT
-- u+2599:
-- 0x8b:
    "11110000",
    "11110000",
    "11110000",
    "11110000",
    "11111111",
    "11111111",
    "11111111",
    "11111111",


-- # [?] QUADRANT UPPER RIGHT AND LOWER LEFT AND LOWER RIGHT
-- u+259f:
-- 0x8c:
    "00001111",
    "00001111",
    "00001111",
    "00001111",
    "11111111",
    "11111111",
    "11111111",
    "11111111",


-- # [?] HORIZONTAL SCAN LINE-1",
-- u+23ba:
-- 0x8d:
    "00000000",
    "00000000",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11111111",


-- # [?] HORIZONTAL SCAN LINE-9
-- u+23bd:
-- 0x8e:
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "00000000",
    "00000000",


-- # [?] QUADRANT UPPER LEFT AND UPPER RIGHT AND LOWER RIGHT
-- u+259c:
-- 0x8f:
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "00001111",
    "00001111",
    "00001111",
    "00001111",


-- # [?] BLACK CLUB SUIT
-- u+2663:
-- 0x90:
    "11111111",
    "11100011",
    "11100011",
    "10001000",
    "10001000",
    "11110111",
    "11100011",
    "11111111",


-- # [?] BOX DRAWINGS LIGHT DOWN AND RIGHT
-- u+250c:
-- 0x91:
    "11111111",
    "11111111",
    "11111111",
    "11100000",
    "11100000",
    "11100111",
    "11100111",
    "11100111",


-- # [?] BOX DRAWINGS LIGHT HORIZONTAL
-- u+2500:
-- 0x92:
    "11111111",
    "11111111",
    "11111111",
    "00000000",
    "00000000",
    "11111111",
    "11111111",
    "11111111",


-- # [?] BOX DRAWINGS LIGHT VERTICAL AND HORIZONTAL
-- u+253c:
-- 0x93:
    "11100111",
    "11100111",
    "11100111",
    "00000000",
    "00000000",
    "11100111",
    "11100111",
    "11100111",


-- # [?] INVERSE BULLET
-- u+25d8:
-- 0x94:
    "11111111",
    "11111111",
    "11000011",
    "10000001",
    "10000001",
    "10000001",
    "11000011",
    "11111111",


-- # [?] UPPER HALF BLOCK
-- u+2580:
-- 0x95:
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "00000000",
    "00000000",
    "00000000",
    "00000000",


-- # [?] LEFT VERTICAL BOX LINE
-- u+23b8:
-- 0x96:
    "00111111",
    "00111111",
    "00111111",
    "00111111",
    "00111111",
    "00111111",
    "00111111",
    "00111111",


-- # [?] BOX DRAWINGS LIGHT DOWN AND HORIZONTAL
-- u+252c:
-- 0x97:
    "11111111",
    "11111111",
    "11111111",
    "00000000",
    "00000000",
    "11100111",
    "11100111",
    "11100111",


-- # [?] BOX DRAWINGS LIGHT UP AND HORIZONTAL
-- u+2534:
-- 0x98:
    "11100111",
    "11100111",
    "11100111",
    "00000000",
    "00000000",
    "11111111",
    "11111111",
    "11111111",


-- # [?] RIGHT HALF BLOCK
-- u+2590:
-- 0x99:
    "00001111",
    "00001111",
    "00001111",
    "00001111",
    "00001111",
    "00001111",
    "00001111",
    "00001111",


-- # [?] BOX DRAWINGS LIGHT UP AND RIGHT
-- u+2514:
-- 0x9a:
    "11100111",
    "11100111",
    "11100111",
    "11100000",
    "11100000",
    "11111111",
    "11111111",
    "11111111",

-- 0x9b:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",

-- 0x9c:
    "11111111",
    "11100111",
    "11000011",
    "10000001",
    "11100111",
    "11100111",
    "11100111",
    "11111111",

-- 0x9d:
    "11111111",
    "11100111",
    "11100111",
    "11100111",
    "10000001",
    "11000011",
    "11100111",
    "11111111",

-- 0x9e:
    "11111111",
    "11100111",
    "11001111",
    "10000001",
    "11001111",
    "11100111",
    "11111111",
    "11111111",

-- 0x9f:
    "11111111",
    "11100111",
    "11110011",
    "10000001",
    "11110011",
    "11100111",
    "11111111",
    "11111111",


-- # [ ] SPACE
-- u+0020:
-- 0xa0:
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11111111",


-- # [!] EXCLAMATION MARK
-- u+0021:
-- 0xa1:
    "11111111",
    "11100111",
    "11100111",
    "11100111",
    "11100111",
    "11111111",
    "11100111",
    "11111111",


-- # ["] QUOTATION MARK
-- u+0022:
-- 0xa2:
    "11111111",
    "10011001",
    "10011001",
    "10011001",
    "11111111",
    "11111111",
    "11111111",
    "11111111",


-- # [-- #] NUMBER SIGN
-- u+0023:
-- 0xa3:
    "11111111",
    "10011001",
    "00000000",
    "10011001",
    "10011001",
    "00000000",
    "10011001",
    "11111111",


-- # [$] DOLLAR SIGN
-- u+0024:
-- 0xa4:
    "11100111",
    "11000001",
    "10011111",
    "11000011",
    "11111001",
    "10000011",
    "11100111",
    "11111111",


-- # [%] PERCENT SIGN
-- u+0025:
-- 0xa5:
    "11111111",
    "10011001",
    "10010011",
    "11100111",
    "11001111",
    "10011001",
    "10111001",
    "11111111",


-- # [&] AMPERSAND
-- u+0026:
-- 0xa6:
    "11100011",
    "11001001",
    "11100011",
    "11000111",
    "10010000",
    "10011001",
    "11000100",
    "11111111",


-- # ['] APOSTROPHE
-- u+0027:
-- 0xa7:
    "11111111",
    "11100111",
    "11100111",
    "11100111",
    "11111111",
    "11111111",
    "11111111",
    "11111111",


-- # [(] LEFT PARENTHESIS
-- u+0028:
-- 0xa8:
    "11111111",
    "11110001",
    "11100011",
    "11100111",
    "11100111",
    "11100011",
    "11110001",
    "11111111",


-- # [)] RIGHT PARENTHESIS
-- u+0029:
-- 0xa9:
    "11111111",
    "10001111",
    "11000111",
    "11100111",
    "11100111",
    "11000111",
    "10001111",
    "11111111",


-- # [*] ASTERISK
-- u+002a:
-- 0xaa:
    "11111111",
    "10011001",
    "11000011",
    "00000000",
    "11000011",
    "10011001",
    "11111111",
    "11111111",


-- # [+] PLUS SIGN
-- u+002b:
-- 0xab:
    "11111111",
    "11100111",
    "11100111",
    "10000001",
    "11100111",
    "11100111",
    "11111111",
    "11111111",


-- # [,] COMMA
-- u+002c:
-- 0xac:
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11100111",
    "11100111",
    "11001111",


-- # [-] HYPHEN-MINUS
-- u+002d:
-- 0xad:
    "11111111",
    "11111111",
    "11111111",
    "10000001",
    "11111111",
    "11111111",
    "11111111",
    "11111111",


-- # [0] FULL STOP
-- u+002e:
-- 0xae:
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11100111",
    "11100111",
    "11111111",


-- # [/] SOLIDUS
-- u+002f:
-- 0xaf:
    "11111111",
    "11111001",
    "11110011",
    "11100111",
    "11001111",
    "10011111",
    "10111111",
    "11111111",


-- # [0] DIGIT ZERO
-- u+0030:
-- 0xb0:
    "11111111",
    "11000011",
    "10011001",
    "10010001",
    "10001001",
    "10011001",
    "11000011",
    "11111111",


-- # [1] DIGIT ONE
-- u+0031:
-- 0xb1:
    "11111111",
    "11100111",
    "11000111",
    "11100111",
    "11100111",
    "11100111",
    "10000001",
    "11111111",


-- # [2] DIGIT TWO
-- u+0032:
-- 0xb2:
    "11111111",
    "11000011",
    "10011001",
    "11110011",
    "11100111",
    "11001111",
    "10000001",
    "11111111",


-- # [3] DIGIT THREE
-- u+0033:
-- 0xb3:
    "11111111",
    "10000001",
    "11110011",
    "11100111",
    "11110011",
    "10011001",
    "11000011",
    "11111111",


-- # [4] DIGIT FOUR
-- u+0034:
-- 0xb4:
    "11111111",
    "11110011",
    "11100011",
    "11000011",
    "10010011",
    "10000001",
    "11110011",
    "11111111",


-- # [5] DIGIT FIVE
-- u+0035:
-- 0xb5:
    "11111111",
    "10000001",
    "10011111",
    "10000011",
    "11111001",
    "10011001",
    "11000011",
    "11111111",


-- # [6] DIGIT SIX
-- u+0036:
-- 0xb6:
    "11111111",
    "11000011",
    "10011111",
    "10000011",
    "10011001",
    "10011001",
    "11000011",
    "11111111",


-- # [7] DIGIT SEVEN
-- u+0037:
-- 0xb7:
    "11111111",
    "10000001",
    "11111001",
    "11110011",
    "11100111",
    "11001111",
    "11001111",
    "11111111",


-- # [8] DIGIT EIGHT
-- u+0038:
-- 0xb8:
    "11111111",
    "11000011",
    "10011001",
    "11000011",
    "10011001",
    "10011001",
    "11000011",
    "11111111",


-- # [9] DIGIT NINE
-- u+0039:
-- 0xb9:
    "11111111",
    "11000011",
    "10011001",
    "11000001",
    "11111001",
    "11110011",
    "11000111",
    "11111111",


-- # [:] COLON
-- u+003a:
-- 0xba:
    "11111111",
    "11111111",
    "11100111",
    "11100111",
    "11111111",
    "11100111",
    "11100111",
    "11111111",


-- # [;] SEMICOLON
-- u+003b:
-- 0xbb:
    "11111111",
    "11111111",
    "11100111",
    "11100111",
    "11111111",
    "11100111",
    "11100111",
    "11001111",


-- # [<] LESS-THAN SIGN
-- u+003c:
-- 0xbc:
    "11111001",
    "11110011",
    "11100111",
    "11001111",
    "11100111",
    "11110011",
    "11111001",
    "11111111",


-- # [=] EQUALS SIGN
-- u+003d:
-- 0xbd:
    "11111111",
    "11111111",
    "10000001",
    "11111111",
    "11111111",
    "10000001",
    "11111111",
    "11111111",


-- # [>] GREATER-THAN SIGN
-- u+003e:
-- 0xbe:
    "10011111",
    "11001111",
    "11100111",
    "11110011",
    "11100111",
    "11001111",
    "10011111",
    "11111111",


-- # [?] QUESTION MARK
-- u+003f:
-- 0xbf:
    "11111111",
    "11000011",
    "10011001",
    "11110011",
    "11100111",
    "11111111",
    "11100111",
    "11111111",


-- # [1] COMMERCIAL AT
-- u+0040:
-- 0xc0:
    "11111111",
    "11000011",
    "10011001",
    "10010001",
    "10010001",
    "10011111",
    "11000001",
    "11111111",


-- # [A] LATIN CAPITAL LETTER A
-- u+0041:
-- 0xc1:
    "11111111",
    "11100111",
    "11000011",
    "10011001",
    "10011001",
    "10000001",
    "10011001",
    "11111111",


-- # [B] LATIN CAPITAL LETTER B
-- u+0042:
-- 0xc2:
    "11111111",
    "10000011",
    "10011001",
    "10000011",
    "10011001",
    "10011001",
    "10000011",
    "11111111",


-- # [C] LATIN CAPITAL LETTER C
-- u+0043:
-- 0xc3:
    "11111111",
    "11000011",
    "10011001",
    "10011111",
    "10011111",
    "10011001",
    "11000011",
    "11111111",


-- # [D] LATIN CAPITAL LETTER D
-- u+0044:
-- 0xc4:
    "11111111",
    "10000111",
    "10010011",
    "10011001",
    "10011001",
    "10010011",
    "10000111",
    "11111111",


-- # [E] LATIN CAPITAL LETTER E
-- u+0045:
-- 0xc5:
    "11111111",
    "10000001",
    "10011111",
    "10000011",
    "10011111",
    "10011111",
    "10000001",
    "11111111",


-- # [F] LATIN CAPITAL LETTER F
-- u+0046:
-- 0xc6:
    "11111111",
    "10000001",
    "10011111",
    "10000011",
    "10011111",
    "10011111",
    "10011111",
    "11111111",


-- # [G] LATIN CAPITAL LETTER G
-- u+0047:
-- 0xc7:
    "11111111",
    "11000001",
    "10011111",
    "10011111",
    "10010001",
    "10011001",
    "11000001",
    "11111111",


-- # [H] LATIN CAPITAL LETTER H
-- u+0048:
-- 0xc8:
    "11111111",
    "10011001",
    "10011001",
    "10000001",
    "10011001",
    "10011001",
    "10011001",
    "11111111",


-- # [I] LATIN CAPITAL LETTER I
-- u+0049:
-- 0xc9:
    "11111111",
    "10000001",
    "11100111",
    "11100111",
    "11100111",
    "11100111",
    "10000001",
    "11111111",


-- # [J] LATIN CAPITAL LETTER J
-- u+004a:
-- 0xca:
    "11111111",
    "11111001",
    "11111001",
    "11111001",
    "11111001",
    "10011001",
    "11000011",
    "11111111",


-- # [K] LATIN CAPITAL LETTER K
-- u+004b:
-- 0xcb:
    "11111111",
    "10011001",
    "10010011",
    "10000111",
    "10000111",
    "10010011",
    "10011001",
    "11111111",


-- # [L] LATIN CAPITAL LETTER L
-- u+004c:
-- 0xcc:
    "11111111",
    "10011111",
    "10011111",
    "10011111",
    "10011111",
    "10011111",
    "10000001",
    "11111111",


-- # [M] LATIN CAPITAL LETTER M
-- u+004d:
-- 0xcd:
    "11111111",
    "10011100",
    "10001000",
    "10000000",
    "10010100",
    "10011100",
    "10011100",
    "11111111",


-- # [N] LATIN CAPITAL LETTER N
-- u+004e:
-- 0xce:
    "11111111",
    "10011001",
    "10001001",
    "10000001",
    "10000001",
    "10010001",
    "10011001",
    "11111111",


-- # [O] LATIN CAPITAL LETTER O
-- u+004f:
-- 0xcf:
    "11111111",
    "11000011",
    "10011001",
    "10011001",
    "10011001",
    "10011001",
    "11000011",
    "11111111",


-- # [P] LATIN CAPITAL LETTER P
-- u+0050:
-- 0xd0:
    "11111111",
    "10000011",
    "10011001",
    "10011001",
    "10000011",
    "10011111",
    "10011111",
    "11111111",


-- # [Q] LATIN CAPITAL LETTER Q
-- u+0051:
-- 0xd1:
    "11111111",
    "11000011",
    "10011001",
    "10011001",
    "10011001",
    "10010011",
    "11001001",
    "11111111",


-- # [R] LATIN CAPITAL LETTER R
-- u+0052:
-- 0xd2:
    "11111111",
    "10000011",
    "10011001",
    "10011001",
    "10000011",
    "10010011",
    "10011001",
    "11111111",


-- # [S] LATIN CAPITAL LETTER S
-- u+0053:
-- 0xd3:
    "11111111",
    "11000011",
    "10011111",
    "11000011",
    "11111001",
    "11111001",
    "11000011",
    "11111111",


-- # [T] LATIN CAPITAL LETTER T
-- u+0054:
-- 0xd4:
    "11111111",
    "10000001",
    "11100111",
    "11100111",
    "11100111",
    "11100111",
    "11100111",
    "11111111",


-- # [U] LATIN CAPITAL LETTER U
-- u+0055:
-- 0xd5:
    "11111111",
    "10011001",
    "10011001",
    "10011001",
    "10011001",
    "10011001",
    "10000001",
    "11111111",


-- # [V] LATIN CAPITAL LETTER V
-- u+0056:
-- 0xd6:
    "11111111",
    "10011001",
    "10011001",
    "10011001",
    "10011001",
    "11000011",
    "11100111",
    "11111111",


-- # [W] LATIN CAPITAL LETTER W
-- u+0057:
-- 0xd7:
    "11111111",
    "10011100",
    "10011100",
    "10010100",
    "10000000",
    "10001000",
    "10011100",
    "11111111",


-- # [X] LATIN CAPITAL LETTER X
-- u+0058:
-- 0xd8:
    "11111111",
    "10011001",
    "10011001",
    "11000011",
    "11000011",
    "10011001",
    "10011001",
    "11111111",


-- # [Y] LATIN CAPITAL LETTER Y
-- u+0059:
-- 0xd9:
    "11111111",
    "10011001",
    "10011001",
    "11000011",
    "11100111",
    "11100111",
    "11100111",
    "11111111",


-- # [Z] LATIN CAPITAL LETTER Z
-- u+005a:
-- 0xda:
    "11111111",
    "10000001",
    "11110011",
    "11100111",
    "11001111",
    "10011111",
    "10000001",
    "11111111",


-- # [[] LEFT SQUARE BRACKET
-- u+005b:
-- 0xdb:
    "11111111",
    "11100001",
    "11100111",
    "11100111",
    "11100111",
    "11100111",
    "11100001",
    "11111111",


-- # [\] REVERSE SOLIDUS
-- u+005c:
-- 0xdc:
    "11111111",
    "10111111",
    "10011111",
    "11001111",
    "11100111",
    "11110011",
    "11111001",
    "11111111",


-- # []] RIGHT SQUARE BRACKET
-- u+005d:
-- 0xdd:
    "11111111",
    "10000111",
    "11100111",
    "11100111",
    "11100111",
    "11100111",
    "10000111",
    "11111111",


-- # [^] CIRCUMFLEX ACCENT
-- u+005e:
-- 0xde:
    "11111111",
    "11110111",
    "11100011",
    "11001001",
    "10011100",
    "11111111",
    "11111111",
    "11111111",


-- # [_] LOW LINE
-- u+005f:
-- 0xdf:
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "11111111",
    "00000000",
    "11111111",


-- # [?] BLACK DIAMOND SUIT
-- u+2666:
-- 0xe0:
    "11111111",
    "11100111",
    "11000011",
    "10000001",
    "10000001",
    "11000011",
    "11100111",
    "11111111",


-- # [a] LATIN SMALL LETTER A
-- u+0061:
-- 0xe1:
    "11111111",
    "11111111",
    "11000011",
    "11111001",
    "11000001",
    "10011001",
    "11000001",
    "11111111",


-- # [b] LATIN SMALL LETTER B
-- u+0062:
-- 0xe2:
    "11111111",
    "10011111",
    "10011111",
    "10000011",
    "10011001",
    "10011001",
    "10000011",
    "11111111",


-- # [c] LATIN SMALL LETTER C
-- u+0063:
-- 0xe3:
    "11111111",
    "11111111",
    "11000011",
    "10011111",
    "10011111",
    "10011111",
    "11000011",
    "11111111",


-- # [d] LATIN SMALL LETTER D
-- u+0064:
-- 0xe4:
    "11111111",
    "11111001",
    "11111001",
    "11000001",
    "10011001",
    "10011001",
    "11000001",
    "11111111",


-- # [e] LATIN SMALL LETTER E
-- u+0065:
-- 0xe5:
    "11111111",
    "11111111",
    "11000011",
    "10011001",
    "10000001",
    "10011111",
    "11000011",
    "11111111",


-- # [f] LATIN SMALL LETTER F
-- u+0066:
-- 0xe6:
    "11111111",
    "11110001",
    "11100111",
    "11000001",
    "11100111",
    "11100111",
    "11100111",
    "11111111",


-- # [g] LATIN SMALL LETTER G
-- u+0067:
-- 0xe7:
    "11111111",
    "11111111",
    "11000001",
    "10011001",
    "10011001",
    "11000001",
    "11111001",
    "10000011",


-- # [h] LATIN SMALL LETTER H
-- u+0068:
-- 0xe8:
    "11111111",
    "10011111",
    "10011111",
    "10000011",
    "10011001",
    "10011001",
    "10011001",
    "11111111",


-- # [i] LATIN SMALL LETTER I
-- u+0069:
-- 0xe9:
    "11111111",
    "11100111",
    "11111111",
    "11000111",
    "11100111",
    "11100111",
    "11000011",
    "11111111",


-- # [j] LATIN SMALL LETTER J
-- u+006a:
-- 0xea:
    "11111111",
    "11111001",
    "11111111",
    "11111001",
    "11111001",
    "11111001",
    "11111001",
    "11000011",


-- # [k] LATIN SMALL LETTER K
-- u+006b:
-- 0xeb:
    "11111111",
    "10011111",
    "10011111",
    "10010011",
    "10000111",
    "10010011",
    "10011001",
    "11111111",


-- # [l] LATIN SMALL LETTER L
-- u+006c:
-- 0xec:
    "11111111",
    "11000111",
    "11100111",
    "11100111",
    "11100111",
    "11100111",
    "11000011",
    "11111111",


-- # [m] LATIN SMALL LETTER M
-- u+006d:
-- 0xed:
    "11111111",
    "11111111",
    "10011001",
    "10000000",
    "10000000",
    "10010100",
    "10011100",
    "11111111",


-- # [n] LATIN SMALL LETTER N
-- u+006e:
-- 0xee:
    "11111111",
    "11111111",
    "10000011",
    "10011001",
    "10011001",
    "10011001",
    "10011001",
    "11111111",


-- # [o] LATIN SMALL LETTER O
-- u+006f:
-- 0xef:
    "11111111",
    "11111111",
    "11000011",
    "10011001",
    "10011001",
    "10011001",
    "11000011",
    "11111111",


-- # [p] LATIN SMALL LETTER P
-- u+0070:
-- 0xf0:
    "11111111",
    "11111111",
    "10000011",
    "10011001",
    "10011001",
    "10000011",
    "10011111",
    "10011111",


-- # [q] LATIN SMALL LETTER Q
-- u+0071:
-- 0xf1:
    "11111111",
    "11111111",
    "11000001",
    "10011001",
    "10011001",
    "11000001",
    "11111001",
    "11111001",


-- # [r] LATIN SMALL LETTER R
-- u+0072:
-- 0xf2:
    "11111111",
    "11111111",
    "10000011",
    "10011001",
    "10011111",
    "10011111",
    "10011111",
    "11111111",


-- # [s] LATIN SMALL LETTER S
-- u+0073:
-- 0xf3:
    "11111111",
    "11111111",
    "11000001",
    "10011111",
    "11000011",
    "11111001",
    "10000011",
    "11111111",


-- # [t] LATIN SMALL LETTER T
-- u+0074:
-- 0xf4:
    "11111111",
    "11100111",
    "10000001",
    "11100111",
    "11100111",
    "11100111",
    "11110001",
    "11111111",


-- # [u] LATIN SMALL LETTER U
-- u+0075:
-- 0xf5:
    "11111111",
    "11111111",
    "10011001",
    "10011001",
    "10011001",
    "10011001",
    "11000001",
    "11111111",


-- # [v] LATIN SMALL LETTER V
-- u+0076:
-- 0xf6:
    "11111111",
    "11111111",
    "10011001",
    "10011001",
    "10011001",
    "11000011",
    "11100111",
    "11111111",


-- # [w] LATIN SMALL LETTER W
-- u+0077:
-- 0xf7:
    "11111111",
    "11111111",
    "10011100",
    "10010100",
    "10000000",
    "11000001",
    "11001001",
    "11111111",


-- # [x] LATIN SMALL LETTER X
-- u+0078:
-- 0xf8:
    "11111111",
    "11111111",
    "10011001",
    "11000011",
    "11100111",
    "11000011",
    "10011001",
    "11111111",


-- # [y] LATIN SMALL LETTER Y
-- u+0079:
-- 0xf9:
    "11111111",
    "11111111",
    "10011001",
    "10011001",
    "10011001",
    "11000001",
    "11110011",
    "10000111",


-- # [z] LATIN SMALL LETTER Z
-- u+007a:
-- 0xfa:
    "11111111",
    "11111111",
    "10000001",
    "11110011",
    "11100111",
    "11001111",
    "10000001",
    "11111111",


-- # [?] BLACK SPADE SUIT
-- u+2660:
-- 0xfb:
    "11111111",
    "11100111",
    "11000011",
    "10000001",
    "10000001",
    "11100111",
    "11000011",
    "11111111",


-- # [|] VERTICAL LINE
-- u+007c:
-- 0xfc:
    "11100111",
    "11100111",
    "11100111",
    "11100111",
    "11100111",
    "11100111",
    "11100111",
    "11100111",

-- 0xfd:
    "11111111",
    "10000001",
    "10000111",
    "10000011",
    "10010001",
    "10011001",
    "11111001",
    "11111111",

-- 0xfe:
    "11110111",
    "11100111",
    "11000111",
    "10000111",
    "11000111",
    "11100111",
    "11110111",
    "11111111",

-- 0xff:
    "11101111",
    "11100111",
    "11100011",
    "11100001",
    "11100011",
    "11100111",
    "11101111",
    "11111111"

	);
begin

    dataOut <= ROM(to_integer(unsigned(addrIn)));
	
end architecture rtl;