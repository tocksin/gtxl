/*
-- @file rom_synth.vhd
-- @brief ROM containing instructions
-- @author Justin Davis
--
    Copyright (C) 2024  Justin Davis

    This program is free software: you can redistribute it and/or modify
    it under the terms of the GNU Affero General Public License as published
    by the Free Software Foundation, either version 3 of the License, or
    (at your option) any later version.

    This program is distributed in the hope that it will be useful,
    but WITHOUT ANY WARRANTY; without even the implied warranty of
    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
    GNU Affero General Public License for more details.

    You should have received a copy of the GNU Affero General Public License
    along with this program.  If not, see <https://www.gnu.org/licenses/>.
------------------------------------------------------------------------------*/
library ieee;           use ieee.std_logic_1164.all;
                        use ieee.numeric_std.all;

library work;           use work.tools_pkg.all;
                        use work.sys_description_pkg.all;

entity rom_synth is 
    port (  iAddr   : in    slv;
            oData   :   out slv(7 downto 0));
end entity rom_synth;

architecture rtl of rom_synth is
    type rom_type is array (0 to (2**iAddr'length)-1) of std_logic_vector(oData'range);
    signal rom : rom_type := ( 
    
 0 =>x"C2",
 1 =>x"00",
 2 =>x"0B",
 3 =>x"00",
 4 =>x"C2",
 5 =>x"01",
 6 =>x"01",
 7 =>x"03",
 8 =>x"60",
 9 =>x"37",
 10 =>x"EC",
 11 =>x"BE",
 12 =>x"FD",
 13 =>x"06",
 14 =>x"10",
 15 =>x"A2",
 16 =>x"18",
 17 =>x"00",
 18 =>x"01",
 19 =>x"08",
 20 =>x"60",
 21 =>x"18",
 22 =>x"F0",
 23 =>x"1A",
 24 =>x"01",
 25 =>x"08",
 26 =>x"80",
 27 =>x"01",
 28 =>x"02",
 29 =>x"00",
 30 =>x"18",
 31 =>x"40",
 32 =>x"C2",
 33 =>x"08",
 34 =>x"60",
 35 =>x"0C",
 36 =>x"F0",
 37 =>x"36",
 38 =>x"01",
 39 =>x"08",
 40 =>x"60",
 41 =>x"06",
 42 =>x"F0",
 43 =>x"40",
 44 =>x"00",
 45 =>x"0E",
 46 =>x"C2",
 47 =>x"06",
 48 =>x"01",
 49 =>x"00",
 50 =>x"15",
 51 =>x"01",
 52 =>x"E3",
 53 =>x"00",
 54 =>x"00",
 55 =>x"8A",
 56 =>x"C2",
 57 =>x"06",
 58 =>x"01",
 59 =>x"00",
 60 =>x"15",
 61 =>x"01",
 62 =>x"E3",
 63 =>x"00",
 64 =>x"C2",
 65 =>x"09",
 66 =>x"00",
 67 =>x"4C",
 68 =>x"C2",
 69 =>x"06",
 70 =>x"01",
 71 =>x"00",
 72 =>x"15",
 73 =>x"01",
 74 =>x"E3",
 75 =>x"00",
 76 =>x"10",
 77 =>x"A2",
 78 =>x"18",
 79 =>x"00",
 80 =>x"00",
 81 =>x"5A",
 82 =>x"C2",
 83 =>x"06",
 84 =>x"01",
 85 =>x"00",
 86 =>x"15",
 87 =>x"01",
 88 =>x"E3",
 89 =>x"00",
 90 =>x"10",
 91 =>x"A2",
 92 =>x"18",
 93 =>x"40",
 94 =>x"01",
 95 =>x"09",
 96 =>x"80",
 97 =>x"01",
 98 =>x"C2",
 99 =>x"09",
 100 =>x"60",
 101 =>x"06",
 102 =>x"02",
 103 =>x"00",
 104 =>x"02",
 105 =>x"00",
 106 =>x"02",
 107 =>x"00",
 108 =>x"02",
 109 =>x"00",
 110 =>x"02",
 111 =>x"00",
 112 =>x"02",
 113 =>x"00",
 114 =>x"02",
 115 =>x"00",
 116 =>x"02",
 117 =>x"00",
 118 =>x"02",
 119 =>x"00",
 120 =>x"02",
 121 =>x"00",
 122 =>x"18",
 123 =>x"00",
 124 =>x"F0",
 125 =>x"84",
 126 =>x"01",
 127 =>x"00",
 128 =>x"15",
 129 =>x"01",
 130 =>x"E3",
 131 =>x"00",
 132 =>x"00",
 133 =>x"0E",
 134 =>x"C2",
 135 =>x"06",
 136 =>x"FC",
 137 =>x"0E",
 138 =>x"10",
 139 =>x"3C",
 140 =>x"18",
 141 =>x"00",
 142 =>x"00",
 143 =>x"8A",
 144 =>x"C2",
 145 =>x"06",
 146 =>x"01",
 147 =>x"08",
 148 =>x"80",
 149 =>x"01",
 150 =>x"C2",
 151 =>x"08",
 152 =>x"60",
 153 =>x"18",
 154 =>x"02",
 155 =>x"00",
 156 =>x"02",
 157 =>x"00",
 158 =>x"02",
 159 =>x"00",
 160 =>x"02",
 161 =>x"00",
 162 =>x"02",
 163 =>x"00",
 164 =>x"02",
 165 =>x"00",
 166 =>x"02",
 167 =>x"00",
 168 =>x"02",
 169 =>x"00",
 170 =>x"18",
 171 =>x"40",
 172 =>x"EC",
 173 =>x"B8",
 174 =>x"00",
 175 =>x"81",
 176 =>x"C2",
 177 =>x"05",
 178 =>x"00",
 179 =>x"E2",
 180 =>x"C2",
 181 =>x"06",
 182 =>x"10",
 183 =>x"F1",
 184 =>x"01",
 185 =>x"00",
 186 =>x"15",
 187 =>x"01",
 188 =>x"E3",
 189 =>x"00",
 190 =>x"00",
 191 =>x"37",
 192 =>x"C2",
 193 =>x"03",
 194 =>x"00",
 195 =>x"E2",
 196 =>x"C2",
 197 =>x"06",
 198 =>x"00",
 199 =>x"52",
 200 =>x"C2",
 201 =>x"07",
 202 =>x"00",
 203 =>x"81",
 204 =>x"C2",
 205 =>x"05",
 206 =>x"62",
 207 =>x"00",
 208 =>x"C2",
 209 =>x"08",
 210 =>x"C2",
 211 =>x"09",
 212 =>x"00",
 213 =>x"00",
 214 =>x"14",
 215 =>x"40",
 216 =>x"C2",
 217 =>x"04",
 218 =>x"01",
 219 =>x"04",
 220 =>x"80",
 221 =>x"01",
 222 =>x"CA",
 223 =>x"00",
 224 =>x"FC",
 225 =>x"D8",
 226 =>x"15",
 227 =>x"05",
 228 =>x"00",
 229 =>x"C0",
 230 =>x"5D",
 231 =>x"00",
 232 =>x"5D",
 233 =>x"00",
 234 =>x"5D",
 235 =>x"00",
 236 =>x"5D",
 237 =>x"00",
 238 =>x"5D",
 239 =>x"00",
 240 =>x"5D",
 241 =>x"00",
 242 =>x"5D",
 243 =>x"00",
 244 =>x"5D",
 245 =>x"00",
 246 =>x"5D",
 247 =>x"00",
 248 =>x"5D",
 249 =>x"00",
 250 =>x"5D",
 251 =>x"00",
 252 =>x"5D",
 253 =>x"00",
 254 =>x"5D",
 255 =>x"00",
 256 =>x"5D",
 257 =>x"00",
 258 =>x"5D",
 259 =>x"00",
 260 =>x"5D",
 261 =>x"00",
 262 =>x"5D",
 263 =>x"00",
 264 =>x"5D",
 265 =>x"00",
 266 =>x"5D",
 267 =>x"00",
 268 =>x"5D",
 269 =>x"00",
 270 =>x"5D",
 271 =>x"00",
 272 =>x"5D",
 273 =>x"00",
 274 =>x"5D",
 275 =>x"00",
 276 =>x"5D",
 277 =>x"00",
 278 =>x"5D",
 279 =>x"00",
 280 =>x"5D",
 281 =>x"00",
 282 =>x"5D",
 283 =>x"00",
 284 =>x"5D",
 285 =>x"00",
 286 =>x"5D",
 287 =>x"00",
 288 =>x"5D",
 289 =>x"00",
 290 =>x"5D",
 291 =>x"00",
 292 =>x"5D",
 293 =>x"00",
 294 =>x"5D",
 295 =>x"00",
 296 =>x"5D",
 297 =>x"00",
 298 =>x"5D",
 299 =>x"00",
 300 =>x"5D",
 301 =>x"00",
 302 =>x"5D",
 303 =>x"00",
 304 =>x"5D",
 305 =>x"00",
 306 =>x"5D",
 307 =>x"00",
 308 =>x"5D",
 309 =>x"00",
 310 =>x"5D",
 311 =>x"00",
 312 =>x"5D",
 313 =>x"00",
 314 =>x"5D",
 315 =>x"00",
 316 =>x"5D",
 317 =>x"00",
 318 =>x"5D",
 319 =>x"00",
 320 =>x"5D",
 321 =>x"00",
 322 =>x"5D",
 323 =>x"00",
 324 =>x"5D",
 325 =>x"00",
 326 =>x"5D",
 327 =>x"00",
 328 =>x"5D",
 329 =>x"00",
 330 =>x"5D",
 331 =>x"00",
 332 =>x"5D",
 333 =>x"00",
 334 =>x"5D",
 335 =>x"00",
 336 =>x"5D",
 337 =>x"00",
 338 =>x"5D",
 339 =>x"00",
 340 =>x"5D",
 341 =>x"00",
 342 =>x"5D",
 343 =>x"00",
 344 =>x"5D",
 345 =>x"00",
 346 =>x"5D",
 347 =>x"00",
 348 =>x"5D",
 349 =>x"00",
 350 =>x"5D",
 351 =>x"00",
 352 =>x"5D",
 353 =>x"00",
 354 =>x"5D",
 355 =>x"00",
 356 =>x"5D",
 357 =>x"00",
 358 =>x"5D",
 359 =>x"00",
 360 =>x"5D",
 361 =>x"00",
 362 =>x"5D",
 363 =>x"00",
 364 =>x"5D",
 365 =>x"00",
 366 =>x"5D",
 367 =>x"00",
 368 =>x"5D",
 369 =>x"00",
 370 =>x"5D",
 371 =>x"00",
 372 =>x"5D",
 373 =>x"00",
 374 =>x"5D",
 375 =>x"00",
 376 =>x"5D",
 377 =>x"00",
 378 =>x"5D",
 379 =>x"00",
 380 =>x"5D",
 381 =>x"00",
 382 =>x"5D",
 383 =>x"00",
 384 =>x"5D",
 385 =>x"00",
 386 =>x"5D",
 387 =>x"00",
 388 =>x"5D",
 389 =>x"00",
 390 =>x"5D",
 391 =>x"00",
 392 =>x"5D",
 393 =>x"00",
 394 =>x"5D",
 395 =>x"00",
 396 =>x"5D",
 397 =>x"00",
 398 =>x"5D",
 399 =>x"00",
 400 =>x"5D",
 401 =>x"00",
 402 =>x"5D",
 403 =>x"00",
 404 =>x"5D",
 405 =>x"00",
 406 =>x"5D",
 407 =>x"00",
 408 =>x"5D",
 409 =>x"00",
 410 =>x"5D",
 411 =>x"00",
 412 =>x"5D",
 413 =>x"00",
 414 =>x"5D",
 415 =>x"00",
 416 =>x"5D",
 417 =>x"00",
 418 =>x"5D",
 419 =>x"00",
 420 =>x"5D",
 421 =>x"00",
 422 =>x"5D",
 423 =>x"00",
 424 =>x"5D",
 425 =>x"00",
 426 =>x"5D",
 427 =>x"00",
 428 =>x"5D",
 429 =>x"00",
 430 =>x"5D",
 431 =>x"00",
 432 =>x"5D",
 433 =>x"00",
 434 =>x"5D",
 435 =>x"00",
 436 =>x"5D",
 437 =>x"00",
 438 =>x"5D",
 439 =>x"00",
 440 =>x"5D",
 441 =>x"00",
 442 =>x"5D",
 443 =>x"00",
 444 =>x"5D",
 445 =>x"00",
 446 =>x"5D",
 447 =>x"00",
 448 =>x"5D",
 449 =>x"00",
 450 =>x"5D",
 451 =>x"00",
 452 =>x"5D",
 453 =>x"00",
 454 =>x"5D",
 455 =>x"00",
 456 =>x"5D",
 457 =>x"00",
 458 =>x"5D",
 459 =>x"00",
 460 =>x"5D",
 461 =>x"00",
 462 =>x"5D",
 463 =>x"00",
 464 =>x"5D",
 465 =>x"00",
 466 =>x"5D",
 467 =>x"00",
 468 =>x"5D",
 469 =>x"00",
 470 =>x"5D",
 471 =>x"00",
 472 =>x"5D",
 473 =>x"00",
 474 =>x"5D",
 475 =>x"00",
 476 =>x"5D",
 477 =>x"00",
 478 =>x"5D",
 479 =>x"00",
 480 =>x"5D",
 481 =>x"00",
 482 =>x"5D",
 483 =>x"00",
 484 =>x"5D",
 485 =>x"00",
 486 =>x"5D",
 487 =>x"00",
 488 =>x"5D",
 489 =>x"00",
 490 =>x"5D",
 491 =>x"00",
 492 =>x"5D",
 493 =>x"00",
 494 =>x"5D",
 495 =>x"00",
 496 =>x"5D",
 497 =>x"00",
 498 =>x"5D",
 499 =>x"00",
 500 =>x"5D",
 501 =>x"00",
 502 =>x"5D",
 503 =>x"00",
 504 =>x"5D",
 505 =>x"00",
 506 =>x"5D",
 507 =>x"00",
 508 =>x"5D",
 509 =>x"00",
 510 =>x"5D",
 511 =>x"00",
 512 =>x"5D",
 513 =>x"00",
 514 =>x"5D",
 515 =>x"00",
 516 =>x"5D",
 517 =>x"00",
 518 =>x"5D",
 519 =>x"00",
 520 =>x"5D",
 521 =>x"00",
 522 =>x"5D",
 523 =>x"00",
 524 =>x"5D",
 525 =>x"00",
 526 =>x"5D",
 527 =>x"00",
 528 =>x"5D",
 529 =>x"00",
 530 =>x"5D",
 531 =>x"00",
 532 =>x"5D",
 533 =>x"00",
 534 =>x"5D",
 535 =>x"00",
 536 =>x"5D",
 537 =>x"00",
 538 =>x"5D",
 539 =>x"00",
 540 =>x"5D",
 541 =>x"00",
 542 =>x"5D",
 543 =>x"00",
 544 =>x"5D",
 545 =>x"00",
 546 =>x"5D",
 547 =>x"00",
 548 =>x"5D",
 549 =>x"00",
 550 =>x"18",
 551 =>x"40",
 552 =>x"00",
 553 =>x"F9",
 554 =>x"6B",
 555 =>x"00",
 556 =>x"EC",
 557 =>x"32",
 558 =>x"14",
 559 =>x"00",
 560 =>x"E0",
 561 =>x"0E",
 562 =>x"02",
 563 =>x"00",
 564 =>x"02",
 565 =>x"00",
 566 =>x"02",
 567 =>x"00",
 568 =>x"02",
 569 =>x"00",
 570 =>x"02",
 571 =>x"00",
 572 =>x"18",
 573 =>x"00",
 574 =>x"02",
 575 =>x"00",
 576 =>x"02",
 577 =>x"00",
 578 =>x"02",
 579 =>x"00",
 580 =>x"02",
 581 =>x"00",
 582 =>x"02",
 583 =>x"00",
 584 =>x"02",
 585 =>x"00",
 586 =>x"02",
 587 =>x"00",
 588 =>x"02",
 589 =>x"00",
 590 =>x"10",
 591 =>x"F0",
 592 =>x"FD",
 593 =>x"07",
 594 =>x"00",
 595 =>x"5E",
 596 =>x"C2",
 597 =>x"07",
 598 =>x"01",
 599 =>x"00",
 600 =>x"15",
 601 =>x"01",
 602 =>x"18",
 603 =>x"40",
 604 =>x"E3",
 605 =>x"00",
 606 =>x"01",
 607 =>x"05",
 608 =>x"80",
 609 =>x"01",
 610 =>x"C2",
 611 =>x"05",
 612 =>x"00",
 613 =>x"52",
 614 =>x"18",
 615 =>x"40",
 616 =>x"C2",
 617 =>x"07",
 618 =>x"01",
 619 =>x"00",
 620 =>x"15",
 621 =>x"01",
 622 =>x"E3",
 623 =>x"00",


    ----------------------------------------------------------
    ------        X Lookup Table                       -------
    ----------------------------------------------------------

    16128 =>x"00", --3F00
    16129 =>x"01", --3F01
    16130 =>x"02", --3F02
    16131 =>x"03", --3F03
    16132 =>x"04", --3F04
    16133 =>x"05", --3F05
    16134 =>x"06", --3F06
    16135 =>x"07", --3F07
    16136 =>x"08", --3F08
    16137 =>x"09", --3F09
    16138 =>x"0A", --3F0A
    16139 =>x"0B", --3F0B
    16140 =>x"0C", --3F0C
    16141 =>x"0D", --3F0D
    16142 =>x"0E", --3F0E
    16143 =>x"0F", --3F0F
    16144 =>x"10", --3F10
    16145 =>x"11", --3F11
    16146 =>x"12", --3F12
    16147 =>x"13", --3F13
    16148 =>x"14", --3F14
    16149 =>x"15", --3F15
    16150 =>x"16", --3F16
    16151 =>x"17", --3F17
    16152 =>x"18", --3F18
    16153 =>x"19", --3F19
    16154 =>x"1A", --3F1A
    16155 =>x"1B", --3F1B
    16156 =>x"1C", --3F1C
    16157 =>x"1D", --3F1D
    16158 =>x"1E", --3F1E
    16159 =>x"1F", --3F1F
    16160 =>x"20", --3F20
    16161 =>x"21", --3F21
    16162 =>x"22", --3F22
    16163 =>x"23", --3F23
    16164 =>x"24", --3F24
    16165 =>x"25", --3F25
    16166 =>x"26", --3F26
    16167 =>x"27", --3F27
    16168 =>x"28", --3F28
    16169 =>x"29", --3F29
    16170 =>x"2A", --3F2A
    16171 =>x"2B", --3F2B
    16172 =>x"2C", --3F2C
    16173 =>x"2D", --3F2D
    16174 =>x"2E", --3F2E
    16175 =>x"2F", --3F2F
    16176 =>x"30", --3F30
    16177 =>x"31", --3F31
    16178 =>x"32", --3F32
    16179 =>x"33", --3F33
    16180 =>x"34", --3F34
    16181 =>x"35", --3F35
    16182 =>x"36", --3F36
    16183 =>x"37", --3F37
    16184 =>x"38", --3F38
    16185 =>x"39", --3F39
    16186 =>x"3A", --3F3A
    16187 =>x"3B", --3F3B
    16188 =>x"3C", --3F3C
    16189 =>x"3D", --3F3D
    16190 =>x"3E", --3F3E
    16191 =>x"3F", --3F3F
    16192 =>x"40", --3F40
    16193 =>x"41", --3F41
    16194 =>x"42", --3F42
    16195 =>x"43", --3F43
    16196 =>x"44", --3F44
    16197 =>x"45", --3F45
    16198 =>x"46", --3F46
    16199 =>x"47", --3F47
    16200 =>x"48", --3F48
    16201 =>x"49", --3F49
    16202 =>x"4A", --3F4A
    16203 =>x"4B", --3F4B
    16204 =>x"4C", --3F4C
    16205 =>x"4D", --3F4D
    16206 =>x"4E", --3F4E
    16207 =>x"4F", --3F4F
    16208 =>x"50", --3F50
    16209 =>x"51", --3F51
    16210 =>x"52", --3F52
    16211 =>x"53", --3F53
    16212 =>x"54", --3F54
    16213 =>x"55", --3F55
    16214 =>x"56", --3F56
    16215 =>x"57", --3F57
    16216 =>x"58", --3F58
    16217 =>x"59", --3F59
    16218 =>x"5A", --3F5A
    16219 =>x"5B", --3F5B
    16220 =>x"5C", --3F5C
    16221 =>x"5D", --3F5D
    16222 =>x"5E", --3F5E
    16223 =>x"5F", --3F5F
    16224 =>x"60", --3F60
    16225 =>x"61", --3F61
    16226 =>x"62", --3F62
    16227 =>x"63", --3F63
    16228 =>x"64", --3F64
    16229 =>x"65", --3F65
    16230 =>x"66", --3F66
    16231 =>x"67", --3F67
    16232 =>x"68", --3F68
    16233 =>x"69", --3F69
    16234 =>x"6A", --3F6A
    16235 =>x"6B", --3F6B
    16236 =>x"6C", --3F6C
    16237 =>x"6D", --3F6D
    16238 =>x"6E", --3F6E
    16239 =>x"6F", --3F6F
    16240 =>x"70", --3F70
    16241 =>x"71", --3F71
    16242 =>x"72", --3F72
    16243 =>x"73", --3F73
    16244 =>x"74", --3F74
    16245 =>x"75", --3F75
    16246 =>x"76", --3F76
    16247 =>x"77", --3F77
    16248 =>x"78", --3F78
    16249 =>x"79", --3F79
    16250 =>x"7A", --3F7A
    16251 =>x"7B", --3F7B
    16252 =>x"7C", --3F7C
    16253 =>x"7D", --3F7D
    16254 =>x"7E", --3F7E
    16255 =>x"7F", --3F7F
    16256 =>x"80", --3F80
    16257 =>x"81", --3F81
    16258 =>x"82", --3F82
    16259 =>x"83", --3F83
    16260 =>x"84", --3F84
    16261 =>x"85", --3F85
    16262 =>x"86", --3F86
    16263 =>x"87", --3F87
    16264 =>x"88", --3F88
    16265 =>x"89", --3F89
    16266 =>x"8A", --3F8A
    16267 =>x"8B", --3F8B
    16268 =>x"8C", --3F8C
    16269 =>x"8D", --3F8D
    16270 =>x"8E", --3F8E
    16271 =>x"8F", --3F8F
    16272 =>x"90", --3F90
    16273 =>x"91", --3F91
    16274 =>x"92", --3F92
    16275 =>x"93", --3F93
    16276 =>x"94", --3F94
    16277 =>x"95", --3F95
    16278 =>x"96", --3F96
    16279 =>x"97", --3F97
    16280 =>x"98", --3F98
    16281 =>x"99", --3F99
    16282 =>x"9A", --3F9A
    16283 =>x"9B", --3F9B
    16284 =>x"9C", --3F9C
    16285 =>x"9D", --3F9D
    16286 =>x"9E", --3F9E
    16287 =>x"9F", --3F9F
    16288 =>x"A0", --3FA0
    16289 =>x"A1", --3FA1
    16290 =>x"A2", --3FA2
    16291 =>x"A3", --3FA3
    16292 =>x"A4", --3FA4
    16293 =>x"A5", --3FA5
    16294 =>x"A6", --3FA6
    16295 =>x"A7", --3FA7
    16296 =>x"A8", --3FA8
    16297 =>x"A9", --3FA9
    16298 =>x"AA", --3FAA
    16299 =>x"AB", --3FAB
    16300 =>x"AC", --3FAC
    16301 =>x"AD", --3FAD
    16302 =>x"AE", --3FAE
    16303 =>x"AF", --3FAF
    16304 =>x"B0", --3FB0
    16305 =>x"B1", --3FB1
    16306 =>x"B2", --3FB2
    16307 =>x"B3", --3FB3
    16308 =>x"B4", --3FB4
    16309 =>x"B5", --3FB5
    16310 =>x"B6", --3FB6
    16311 =>x"B7", --3FB7
    16312 =>x"B8", --3FB8
    16313 =>x"B9", --3FB9
    16314 =>x"BA", --3FBA
    16315 =>x"BB", --3FBB
    16316 =>x"BC", --3FBC
    16317 =>x"BD", --3FBD
    16318 =>x"BE", --3FBE
    16319 =>x"BF", --3FBF
    16320 =>x"C0", --3FC0
    16321 =>x"C1", --3FC1
    16322 =>x"C2", --3FC2
    16323 =>x"C3", --3FC3
    16324 =>x"C4", --3FC4
    16325 =>x"C5", --3FC5
    16326 =>x"C6", --3FC6
    16327 =>x"C7", --3FC7
    16328 =>x"C8", --3FC8
    16329 =>x"C9", --3FC9
    16330 =>x"CA", --3FCA
    16331 =>x"CB", --3FCB
    16332 =>x"CC", --3FCC
    16333 =>x"CD", --3FCD
    16334 =>x"CE", --3FCE
    16335 =>x"CF", --3FCF
    16336 =>x"D0", --3FD0
    16337 =>x"D1", --3FD1
    16338 =>x"D2", --3FD2
    16339 =>x"D3", --3FD3
    16340 =>x"D4", --3FD4
    16341 =>x"D5", --3FD5
    16342 =>x"D6", --3FD6
    16343 =>x"D7", --3FD7
    16344 =>x"D8", --3FD8
    16345 =>x"D9", --3FD9
    16346 =>x"DA", --3FDA
    16347 =>x"DB", --3FDB
    16348 =>x"DC", --3FDC
    16349 =>x"DD", --3FDD
    16350 =>x"DE", --3FDE
    16351 =>x"DF", --3FDF
    16352 =>x"E0", --3FE0
    16353 =>x"E1", --3FE1
    16354 =>x"E2", --3FE2
    16355 =>x"E3", --3FE3
    16356 =>x"E4", --3FE4
    16357 =>x"E5", --3FE5
    16358 =>x"E6", --3FE6
    16359 =>x"E7", --3FE7
    16360 =>x"E8", --3FE8
    16361 =>x"E9", --3FE9
    16362 =>x"EA", --3FEA
    16363 =>x"EB", --3FEB
    16364 =>x"EC", --3FEC
    16365 =>x"ED", --3FED
    16366 =>x"EE", --3FEE
    16367 =>x"EF", --3FEF
    16368 =>x"F0", --3FF0
    16369 =>x"F1", --3FF1
    16370 =>x"F2", --3FF2
    16371 =>x"F3", --3FF3
    16372 =>x"F4", --3FF4
    16373 =>x"F5", --3FF5
    16374 =>x"F6", --3FF6
    16375 =>x"F7", --3FF7
    16376 =>x"F8", --3FF8
    16377 =>x"F9", --3FF9
    16378 =>x"FA", --3FFA
    16379 =>x"FB", --3FFB
    16380 =>x"FC", --3FFC
    16381 =>x"FD", --3FFD
    16382 =>x"FE", --3FFE
    16383 =>x"FF", --3FFF


    others => (others=>'0')
    );

begin
       oData <= rom(to_integer(unsigned(iAddr)));
end rtl;
