-- @file rom_font.vhd
-- @brief ROM containing character font
-- @author Justin Davis
--
-- $Revision: -
-- $Date: 06/22/2023
-- $LastEditedBy: Justin Davis
--
-- Developed by 2023 Southwest Research Institute
-------------------------------------------------------------------------------
-- Font data taken from: https://github.com/robhagemans/hoard-of-bitfonts/blob/master/commodore/pet/pet.yaff

library ieee;           use ieee.std_logic_1164.all;
                        use ieee.numeric_std.all;

library work;           use work.tools_pkg.all;
                        use work.sys_description_pkg.all;

entity rom_font is
    port ( addrIn   : in    slv(10 downto 0) ;
           dataOut  :   out slv(7 downto 0));
end entity rom_font;

architecture rtl of rom_font is
   
    type rom_type is array (0 to (2**addrIn'length)-1) of std_logic_vector(dataOut'range);

    -- ROM definition
    signal rom : rom_type := ( 

-- # [1] COMMERCIAL AT
-- 0x00:
-- u+0040:
    "00011100",
    "00100010",
    "01001010",
    "01010110",
    "01001100",
    "00100000",
    "00011110",
    "00000000",


-- # [A] LATIN CAPITAL LETTER A
-- 0x01:
-- u+0041:
    "00011000",
    "00100100",
    "01000010",
    "01111110",
    "01000010",
    "01000010",
    "01000010",
    "00000000",


-- # [B] LATIN CAPITAL LETTER B
-- 0x02:
-- u+0042:
    "01111100",
    "00100010",
    "00100010",
    "00111100",
    "00100010",
    "00100010",
    "01111100",
    "00000000",


-- # [C] LATIN CAPITAL LETTER C
-- 0x03:
-- u+0043:
    "00011100",
    "00100010",
    "01000000",
    "01000000",
    "01000000",
    "00100010",
    "00011100",
    "00000000",


-- # [D] LATIN CAPITAL LETTER D
-- 0x04:
-- u+0044:
    "01111000",
    "00100100",
    "00100010",
    "00100010",
    "00100010",
    "00100100",
    "01111000",
    "00000000",


-- # [E] LATIN CAPITAL LETTER E
-- 0x05:
-- u+0045:
    "01111110",
    "01000000",
    "01000000",
    "01111000",
    "01000000",
    "01000000",
    "01111110",
    "00000000",


-- # [F] LATIN CAPITAL LETTER F
-- 0x06:
-- u+0046:
    "01111110",
    "01000000",
    "01000000",
    "01111000",
    "01000000",
    "01000000",
    "01000000",
    "00000000",


-- # [G] LATIN CAPITAL LETTER G
-- 0x07:
-- u+0047:
    "00011100",
    "00100010",
    "01000000",
    "01001110",
    "01000010",
    "00100010",
    "00011100",
    "00000000",


-- # [H] LATIN CAPITAL LETTER H
-- 0x08:
-- u+0048:
    "01000010",
    "01000010",
    "01000010",
    "01111110",
    "01000010",
    "01000010",
    "01000010",
    "00000000",


-- # [I] LATIN CAPITAL LETTER I
-- 0x09:
-- u+0049:
    "00011100",
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00011100",
    "00000000",


-- # [J] LATIN CAPITAL LETTER J
-- 0x0a:
-- u+004a:
    "00001110",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "01000100",
    "00111000",
    "00000000",


-- # [K] LATIN CAPITAL LETTER K
-- 0x0b:
-- u+004b:
    "01000010",
    "01000100",
    "01001000",
    "01110000",
    "01001000",
    "01000100",
    "01000010",
    "00000000",


-- # [L] LATIN CAPITAL LETTER L
-- 0x0c:
-- u+004c:
    "01000000",
    "01000000",
    "01000000",
    "01000000",
    "01000000",
    "01000000",
    "01111110",
    "00000000",


-- # [M] LATIN CAPITAL LETTER M
-- 0x0d:
-- u+004d:
    "01000010",
    "01100110",
    "01011010",
    "01011010",
    "01000010",
    "01000010",
    "01000010",
    "00000000",


-- # [N] LATIN CAPITAL LETTER N
-- 0x0e:
-- u+004e:
    "01000010",
    "01100010",
    "01010010",
    "01001010",
    "01000110",
    "01000010",
    "01000010",
    "00000000",


-- # [O] LATIN CAPITAL LETTER O
-- 0x0f:
-- u+004f:
    "00011000",
    "00100100",
    "01000010",
    "01000010",
    "01000010",
    "00100100",
    "00011000",
    "00000000",


-- # [P] LATIN CAPITAL LETTER P
-- 0x10:
-- u+0050:
    "01111100",
    "01000010",
    "01000010",
    "01111100",
    "01000000",
    "01000000",
    "01000000",
    "00000000",


-- # [Q] LATIN CAPITAL LETTER Q
-- 0x11:
-- u+0051:
    "00011000",
    "00100100",
    "01000010",
    "01000010",
    "01001010",
    "00100100",
    "00011010",
    "00000000",


-- # [R] LATIN CAPITAL LETTER R
-- 0x12:
-- u+0052:
    "01111100",
    "01000010",
    "01000010",
    "01111100",
    "01001000",
    "01000100",
    "01000010",
    "00000000",


-- # [S] LATIN CAPITAL LETTER S
-- 0x13:
-- u+0053:
    "00111100",
    "01000010",
    "01000000",
    "00111100",
    "00000010",
    "01000010",
    "00111100",
    "00000000",


-- # [T] LATIN CAPITAL LETTER T
-- 0x14:
-- u+0054:
    "00111110",
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00000000",


-- # [U] LATIN CAPITAL LETTER U
-- 0x15:
-- u+0055:
    "01000010",
    "01000010",
    "01000010",
    "01000010",
    "01000010",
    "01000010",
    "00111100",
    "00000000",


-- # [V] LATIN CAPITAL LETTER V
-- 0x16:
-- u+0056:
    "01000010",
    "01000010",
    "01000010",
    "00100100",
    "00100100",
    "00011000",
    "00011000",
    "00000000",


-- # [W] LATIN CAPITAL LETTER W
-- 0x17:
-- u+0057:
    "01000010",
    "01000010",
    "01000010",
    "01011010",
    "01011010",
    "01100110",
    "01000010",
    "00000000",


-- # [X] LATIN CAPITAL LETTER X
-- 0x18:
-- u+0058:
    "01000010",
    "01000010",
    "00100100",
    "00011000",
    "00100100",
    "01000010",
    "01000010",
    "00000000",


-- # [Y] LATIN CAPITAL LETTER Y
-- 0x19:
-- u+0059:
    "00100010",
    "00100010",
    "00100010",
    "00011100",
    "00001000",
    "00001000",
    "00001000",
    "00000000",


-- # [Z] LATIN CAPITAL LETTER Z
-- 0x1a:
-- u+005a:
    "01111110",
    "00000010",
    "00000100",
    "00011000",
    "00100000",
    "01000000",
    "01111110",
    "00000000",


-- # [[] LEFT SQUARE BRACKET
-- 0x1b:
-- u+005b:
    "00111100",
    "00100000",
    "00100000",
    "00100000",
    "00100000",
    "00100000",
    "00111100",
    "00000000",


-- # [\] REVERSE SOLIDUS
-- 0x1c:
-- u+005c:
    "00000000",
    "01000000",
    "00100000",
    "00010000",
    "00001000",
    "00000100",
    "00000010",
    "00000000",


-- # []] RIGHT SQUARE BRACKET
-- 0x1d:
-- u+005d:
    "00111100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00111100",
    "00000000",


-- # [↑] UPWARDS ARROW
-- 0x1e:
-- u+2191:
    "00000000",
    "00001000",
    "00011100",
    "00101010",
    "00001000",
    "00001000",
    "00001000",
    "00001000",


-- # [←] LEFTWARDS ARROW
-- 0x1f:
-- u+2190:
    "00000000",
    "00000000",
    "00010000",
    "00100000",
    "01111111",
    "00100000",
    "00010000",
    "00000000",


-- # [ ] SPACE
-- 0x20:
-- u+0020:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",


-- # [!] EXCLAMATION MARK
-- 0x21:
-- u+0021:
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00000000",
    "00000000",
    "00001000",
    "00000000",


-- # ["] QUOTATION MARK
-- 0x22:
-- u+0022:
    "00100100",
    "00100100",
    "00100100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",


-- # [-- #] NUMBER SIGN
-- 0x23:
-- u+0023:
    "00100100",
    "00100100",
    "01111110",
    "00100100",
    "01111110",
    "00100100",
    "00100100",
    "00000000",


-- # [$] DOLLAR SIGN
-- 0x24:
-- u+0024:
    "00001000",
    "00011110",
    "00101000",
    "00011100",
    "00001010",
    "00111100",
    "00001000",
    "00000000",


-- # [%] PERCENT SIGN
-- 0x25:
-- u+0025:
    "00000000",
    "01100010",
    "01100100",
    "00001000",
    "00010000",
    "00100110",
    "01000110",
    "00000000",


-- # [&] AMPERSAND
-- 0x26:
-- u+0026:
    "00110000",
    "01001000",
    "01001000",
    "00110000",
    "01001010",
    "01000100",
    "00111010",
    "00000000",


-- # ['] APOSTROPHE
-- 0x27:
-- u+0027:
    "00000100",
    "00001000",
    "00010000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",


-- # [(] LEFT PARENTHESIS
-- 0x28:
-- u+0028:
    "00000100",
    "00001000",
    "00010000",
    "00010000",
    "00010000",
    "00001000",
    "00000100",
    "00000000",


-- # [)] RIGHT PARENTHESIS
-- 0x29:
-- u+0029:
    "00100000",
    "00010000",
    "00001000",
    "00001000",
    "00001000",
    "00010000",
    "00100000",
    "00000000",


-- # [*] ASTERISK
-- 0x2a:
-- u+002a:
    "00001000",
    "00101010",
    "00011100",
    "00111110",
    "00011100",
    "00101010",
    "00001000",
    "00000000",


-- # [+] PLUS SIGN
-- 0x2b:
-- u+002b:
    "00000000",
    "00001000",
    "00001000",
    "00111110",
    "00001000",
    "00001000",
    "00000000",
    "00000000",


-- # [,] COMMA
-- 0x2c:
-- u+002c:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00001000",
    "00001000",
    "00010000",


-- # [-] HYPHEN-MINUS
-- 0x2d:
-- u+002d:
    "00000000",
    "00000000",
    "00000000",
    "01111110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",


-- # [0] FULL STOP
-- 0x2e:
-- u+002e:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011000",
    "00011000",
    "00000000",


-- # [/] SOLIDUS
-- 0x2f:
-- u+002f:
    "00000000",
    "00000010",
    "00000100",
    "00001000",
    "00010000",
    "00100000",
    "01000000",
    "00000000",


-- # [0] DIGIT ZERO
-- 0x30:
-- u+0030:
    "00111100",
    "01000010",
    "01000110",
    "01011010",
    "01100010",
    "01000010",
    "00111100",
    "00000000",


-- # [1] DIGIT ONE
-- 0x31:
-- u+0031:
    "00001000",
    "00011000",
    "00101000",
    "00001000",
    "00001000",
    "00001000",
    "00111110",
    "00000000",


-- # [2] DIGIT TWO
-- 0x32:
-- u+0032:
    "00111100",
    "01000010",
    "00000010",
    "00001100",
    "00110000",
    "01000000",
    "01111110",
    "00000000",


-- # [3] DIGIT THREE
-- 0x33:
-- u+0033:
    "00111100",
    "01000010",
    "00000010",
    "00011100",
    "00000010",
    "01000010",
    "00111100",
    "00000000",


-- # [4] DIGIT FOUR
-- 0x34:
-- u+0034:
    "00000100",
    "00001100",
    "00010100",
    "00100100",
    "01111110",
    "00000100",
    "00000100",
    "00000000",


-- # [5] DIGIT FIVE
-- 0x35:
-- u+0035:
    "01111110",
    "01000000",
    "01111000",
    "00000100",
    "00000010",
    "01000100",
    "00111000",
    "00000000",


-- # [6] DIGIT SIX
-- 0x36:
-- u+0036:
    "00011100",
    "00100000",
    "01000000",
    "01111100",
    "01000010",
    "01000010",
    "00111100",
    "00000000",


-- # [7] DIGIT SEVEN
-- 0x37:
-- u+0037:
    "01111110",
    "01000010",
    "00000100",
    "00001000",
    "00010000",
    "00010000",
    "00010000",
    "00000000",


-- # [8] DIGIT EIGHT
-- 0x38:
-- u+0038:
    "00111100",
    "01000010",
    "01000010",
    "00111100",
    "01000010",
    "01000010",
    "00111100",
    "00000000",


-- # [9] DIGIT NINE
-- 0x39:
-- u+0039:
    "00111100",
    "01000010",
    "01000010",
    "00111110",
    "00000010",
    "00000100",
    "00111000",
    "00000000",


-- # [:] COLON
-- 0x3a:
-- u+003a:
    "00000000",
    "00000000",
    "00001000",
    "00000000",
    "00000000",
    "00001000",
    "00000000",
    "00000000",


-- # [;] SEMICOLON
-- 0x3b:
-- u+003b:
    "00000000",
    "00000000",
    "00001000",
    "00000000",
    "00000000",
    "00001000",
    "00001000",
    "00010000",


-- # [<] LESS-THAN SIGN
-- 0x3c:
-- u+003c:
    "00001110",
    "00011000",
    "00110000",
    "01100000",
    "00110000",
    "00011000",
    "00001110",
    "00000000",


-- # [=] EQUALS SIGN
-- 0x3d:
-- u+003d:
    "00000000",
    "00000000",
    "01111110",
    "00000000",
    "01111110",
    "00000000",
    "00000000",
    "00000000",


-- # [>] GREATER-THAN SIGN
-- 0x3e:
-- u+003e:
    "01110000",
    "00011000",
    "00001100",
    "00000110",
    "00001100",
    "00011000",
    "01110000",
    "00000000",


-- # [?] QUESTION MARK
-- 0x3f:
-- u+003f:
    "00111100",
    "01000010",
    "00000010",
    "00001100",
    "00010000",
    "00000000",
    "00010000",
    "00000000",


-- # [─] BOX DRAWINGS LIGHT HORIZONTAL
-- 0x40:
-- u+2500:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111111",
    "00000000",
    "00000000",
    "00000000",


-- # [♠] BLACK SPADE SUIT
-- 0x41:
-- u+2660:
    "00001000",
    "00011100",
    "00111110",
    "01111111",
    "01111111",
    "00011100",
    "00111110",
    "00000000",


-- # [🭲] VERTICAL ONE EIGHTH BLOCK-4
-- 0x42:
-- u+1fb72:
    "00010000",
    "00010000",
    "00010000",
    "00010000",
    "00010000",
    "00010000",
    "00010000",
    "00010000",


-- # [🭸] HORIZONTAL ONE EIGHTH BLOCK-4
-- 0x43:
-- u+1fb78:
    "00000000",
    "00000000",
    "00000000",
    "11111111",
    "00000000",
    "00000000",
    "00000000",
    "00000000",


-- # [🭷] HORIZONTAL ONE EIGHTH BLOCK-3
-- 0x44:
-- u+1fb77:
    "00000000",
    "00000000",
    "11111111",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",


-- # [🭶] HORIZONTAL ONE EIGHTH BLOCK-2
-- 0x45:
-- u+1fb76:
    "00000000",
    "11111111",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",


-- # [🭺] HORIZONTAL ONE EIGHTH BLOCK-6
-- 0x46:
-- u+1fb7a:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111111",
    "00000000",
    "00000000",


-- # [🭱] VERTICAL ONE EIGHTH BLOCK-3
-- 0x47:
-- u+1fb71:
    "00100000",
    "00100000",
    "00100000",
    "00100000",
    "00100000",
    "00100000",
    "00100000",
    "00100000",


-- # [🭴] VERTICAL ONE EIGHTH BLOCK-6
-- 0x48:
-- u+1fb74:
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",


-- # [╮] BOX DRAWINGS LIGHT ARC DOWN AND LEFT
-- 0x49:
-- u+256e:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11100000",
    "00010000",
    "00001000",
    "00001000",


-- # [╰] BOX DRAWINGS LIGHT ARC UP AND RIGHT
-- 0x4a:
-- u+2570:
    "00001000",
    "00001000",
    "00001000",
    "00000100",
    "00000011",
    "00000000",
    "00000000",
    "00000000",


-- # [╯] BOX DRAWINGS LIGHT ARC UP AND LEFT
-- 0x4b:
-- u+256f:
    "00001000",
    "00001000",
    "00001000",
    "00010000",
    "11100000",
    "00000000",
    "00000000",
    "00000000",


-- # [🭼] LEFT AND LOWER ONE EIGHTH BLOCK
-- 0x4c:
-- u+1fb7c:
    "10000000",
    "10000000",
    "10000000",
    "10000000",
    "10000000",
    "10000000",
    "10000000",
    "11111111",


-- # [╲] BOX DRAWINGS LIGHT DIAGONAL UPPER LEFT TO LOWER RIGHT
-- 0x4d:
-- u+2572:
    "10000000",
    "01000000",
    "00100000",
    "00010000",
    "00001000",
    "00000100",
    "00000010",
    "00000001",


-- # [╱] BOX DRAWINGS LIGHT DIAGONAL UPPER RIGHT TO LOWER LEFT
-- 0x4e:
-- u+2571:
    "00000001",
    "00000010",
    "00000100",
    "00001000",
    "00010000",
    "00100000",
    "01000000",
    "10000000",


-- # [🭽] LEFT AND UPPER ONE EIGHTH BLOCK
-- 0x4f:
-- u+1fb7d:
    "11111111",
    "10000000",
    "10000000",
    "10000000",
    "10000000",
    "10000000",
    "10000000",
    "10000000",


-- # [🭾] RIGHT AND UPPER ONE EIGHTH BLOCK
-- 0x50:
-- u+1fb7e:
    "11111111",
    "00000001",
    "00000001",
    "00000001",
    "00000001",
    "00000001",
    "00000001",
    "00000001",


-- # [•] BULLET
-- 0x51:
-- u+2022:
    "00000000",
    "00111100",
    "01111110",
    "01111110",
    "01111110",
    "01111110",
    "00111100",
    "00000000",


-- # [🭻] HORIZONTAL ONE EIGHTH BLOCK-7
-- 0x52:
-- u+1fb7b:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111111",
    "00000000",


-- # [♥] BLACK HEART SUIT
-- 0x53:
-- u+2665:
    "00110110",
    "01111111",
    "01111111",
    "01111111",
    "00111110",
    "00011100",
    "00001000",
    "00000000",


-- # [🭰] VERTICAL ONE EIGHTH BLOCK-2
-- 0x54:
-- u+1fb70:
    "01000000",
    "01000000",
    "01000000",
    "01000000",
    "01000000",
    "01000000",
    "01000000",
    "01000000",


-- # [╭] BOX DRAWINGS LIGHT ARC DOWN AND RIGHT
-- 0x55:
-- u+256d:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000011",
    "00000100",
    "00001000",
    "00001000",


-- # [╳] BOX DRAWINGS LIGHT DIAGONAL CROSS
-- 0x56:
-- u+2573:
    "10000001",
    "01000010",
    "00100100",
    "00011000",
    "00011000",
    "00100100",
    "01000010",
    "10000001",


-- # [○] WHITE CIRCLE
-- 0x57:
-- u+25cb:
    "00000000",
    "00111100",
    "01000010",
    "01000010",
    "01000010",
    "01000010",
    "00111100",
    "00000000",


-- # [♣] BLACK CLUB SUIT
-- 0x58:
-- u+2663:
    "00001000",
    "00011100",
    "00101010",
    "01110111",
    "00101010",
    "00001000",
    "00001000",
    "00000000",


-- # [🭵] VERTICAL ONE EIGHTH BLOCK-7
-- 0x59:
-- u+1fb75:
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",
    "00000010",


-- # [♦] BLACK DIAMOND SUIT
-- 0x5a:
-- u+2666:
    "00001000",
    "00011100",
    "00111110",
    "01111111",
    "00111110",
    "00011100",
    "00001000",
    "00000000",


-- # [┼] BOX DRAWINGS LIGHT VERTICAL AND HORIZONTAL
-- 0x5b:
-- u+253c:
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "11111111",
    "00001000",
    "00001000",
    "00001000",


-- # [🮌] LEFT HALF MEDIUM SHADE
-- 0x5c:
-- u+1fb8c:
    "10100000",
    "01010000",
    "10100000",
    "01010000",
    "10100000",
    "01010000",
    "10100000",
    "01010000",


-- # [│] BOX DRAWINGS LIGHT VERTICAL
-- 0x5d:
-- u+2502:
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00001000",


-- # [π] GREEK SMALL LETTER PI
-- 0x5e:
-- u+03c0:
    "00000000",
    "00000000",
    "00000001",
    "00111110",
    "01010100",
    "00010100",
    "00010100",
    "00000000",


-- # [◥] BLACK UPPER RIGHT TRIANGLE
-- 0x5f:
-- u+25e5:
    "11111111",
    "01111111",
    "00111111",
    "00011111",
    "00001111",
    "00000111",
    "00000011",
    "00000001",


-- # [ ] NO-BREAK SPACE
-- 0x60:
-- u+00a0:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",


-- # [▌] LEFT HALF BLOCK
-- 0x61:
-- u+258c:
    "11110000",
    "11110000",
    "11110000",
    "11110000",
    "11110000",
    "11110000",
    "11110000",
    "11110000",


-- # [▄] LOWER HALF BLOCK
-- 0x62:
-- u+2584:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111111",
    "11111111",
    "11111111",
    "11111111",


-- # [▔] UPPER ONE EIGHTH BLOCK
-- 0x63:
-- u+2594:
    "11111111",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",


-- # [▁] LOWER ONE EIGHTH BLOCK
-- 0x64:
-- u+2581:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111111",


-- # [▏] LEFT ONE EIGHTH BLOCK
-- 0x65:
-- u+258f:
    "10000000",
    "10000000",
    "10000000",
    "10000000",
    "10000000",
    "10000000",
    "10000000",
    "10000000",


-- # [▒] MEDIUM SHADE
-- 0x66:
-- u+2592:
    "10101010",
    "01010101",
    "10101010",
    "01010101",
    "10101010",
    "01010101",
    "10101010",
    "01010101",


-- # [▕] RIGHT ONE EIGHTH BLOCK
-- 0x67:
-- u+2595:
    "00000001",
    "00000001",
    "00000001",
    "00000001",
    "00000001",
    "00000001",
    "00000001",
    "00000001",


-- # [🮏] LOWER HALF MEDIUM SHADE
-- 0x68:
-- u+1fb8f:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "10101010",
    "01010101",
    "10101010",
    "01010101",


-- # [◤] BLACK UPPER LEFT TRIANGLE
-- 0x69:
-- u+25e4:
    "11111111",
    "11111110",
    "11111100",
    "11111000",
    "11110000",
    "11100000",
    "11000000",
    "10000000",


-- # [🮇] RIGHT ONE QUARTER BLOCK
-- 0x6a:
-- u+1fb87:
    "00000011",
    "00000011",
    "00000011",
    "00000011",
    "00000011",
    "00000011",
    "00000011",
    "00000011",


-- # [├] BOX DRAWINGS LIGHT VERTICAL AND RIGHT
-- 0x6b:
-- u+251c:
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00001111",
    "00001000",
    "00001000",
    "00001000",


-- # [▗] QUADRANT LOWER RIGHT
-- 0x6c:
-- u+2597:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00001111",
    "00001111",
    "00001111",
    "00001111",


-- # [└] BOX DRAWINGS LIGHT UP AND RIGHT
-- 0x6d:
-- u+2514:
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00001111",
    "00000000",
    "00000000",
    "00000000",


-- # [┐] BOX DRAWINGS LIGHT DOWN AND LEFT
-- 0x6e:
-- u+2510:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111000",
    "00001000",
    "00001000",
    "00001000",


-- # [▂] LOWER ONE QUARTER BLOCK
-- 0x6f:
-- u+2582:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111111",
    "11111111",


-- # [┌] BOX DRAWINGS LIGHT DOWN AND RIGHT
-- 0x70:
-- u+250c:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00001111",
    "00001000",
    "00001000",
    "00001000",


-- # [┴] BOX DRAWINGS LIGHT UP AND HORIZONTAL
-- 0x71:
-- u+2534:
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "11111111",
    "00000000",
    "00000000",
    "00000000",


-- # [┬] BOX DRAWINGS LIGHT DOWN AND HORIZONTAL
-- 0x72:
-- u+252c:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111111",
    "00001000",
    "00001000",
    "00001000",


-- # [┤] BOX DRAWINGS LIGHT VERTICAL AND LEFT
-- 0x73:
-- u+2524:
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "11111000",
    "00001000",
    "00001000",
    "00001000",


-- # [▎] LEFT ONE QUARTER BLOCK
-- 0x74:
-- u+258e:
    "11000000",
    "11000000",
    "11000000",
    "11000000",
    "11000000",
    "11000000",
    "11000000",
    "11000000",


-- # [▍] LEFT THREE EIGHTHS BLOCK
-- 0x75:
-- u+258d:
    "11100000",
    "11100000",
    "11100000",
    "11100000",
    "11100000",
    "11100000",
    "11100000",
    "11100000",


-- # [🮈] RIGHT THREE EIGHTHS BLOCK
-- 0x76:
-- u+1fb88:
    "00000111",
    "00000111",
    "00000111",
    "00000111",
    "00000111",
    "00000111",
    "00000111",
    "00000111",


-- # [🮂] UPPER ONE QUARTER BLOCK
-- 0x77:
-- u+1fb82:
    "11111111",
    "11111111",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",


-- # [🮃] UPPER THREE EIGHTHS BLOCK
-- 0x78:
-- u+1fb83:
    "11111111",
    "11111111",
    "11111111",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",


-- # [▃] LOWER THREE EIGHTHS BLOCK
-- 0x79:
-- u+2583:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111111",
    "11111111",
    "11111111",


-- # [🭿] RIGHT AND LOWER ONE EIGHTH BLOCK
-- 0x7a:
-- u+1fb7f:
    "00000001",
    "00000001",
    "00000001",
    "00000001",
    "00000001",
    "00000001",
    "00000001",
    "11111111",


-- # [▖] QUADRANT LOWER LEFT
-- 0x7b:
-- u+2596:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11110000",
    "11110000",
    "11110000",
    "11110000",


-- # [▝] QUADRANT UPPER RIGHT
-- 0x7c:
-- u+259d:
    "00001111",
    "00001111",
    "00001111",
    "00001111",
    "00000000",
    "00000000",
    "00000000",
    "00000000",


-- # [┘] BOX DRAWINGS LIGHT UP AND LEFT
-- 0x7d:
-- u+2518:
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "11111000",
    "00000000",
    "00000000",
    "00000000",


-- # [▘] QUADRANT UPPER LEFT
-- 0x7e:
-- u+2598:
    "11110000",
    "11110000",
    "11110000",
    "11110000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",


-- # [▚] QUADRANT UPPER LEFT AND LOWER RIGHT
-- 0x7f:
-- u+259a:
    "11110000",
    "11110000",
    "11110000",
    "11110000",
    "00001111",
    "00001111",
    "00001111",
    "00001111",


-- # [1] COMMERCIAL AT
-- 0x80:
-- u+0040:
    "00011100",
    "00100010",
    "01001010",
    "01010110",
    "01001100",
    "00100000",
    "00011110",
    "00000000",


-- # [a] LATIN SMALL LETTER A
-- 0x81:
-- u+0061:
    "00000000",
    "00000000",
    "00111000",
    "00000100",
    "00111100",
    "01000100",
    "00111010",
    "00000000",


-- # [b] LATIN SMALL LETTER B
-- 0x82:
-- u+0062:
    "01000000",
    "01000000",
    "01011100",
    "01100010",
    "01000010",
    "01100010",
    "01011100",
    "00000000",


-- # [c] LATIN SMALL LETTER C
-- 0x83:
-- u+0063:
    "00000000",
    "00000000",
    "00111100",
    "01000010",
    "01000000",
    "01000010",
    "00111100",
    "00000000",


-- # [d] LATIN SMALL LETTER D
-- 0x84:
-- u+0064:
    "00000010",
    "00000010",
    "00111010",
    "01000110",
    "01000010",
    "01000110",
    "00111010",
    "00000000",


-- # [e] LATIN SMALL LETTER E
-- 0x85:
-- u+0065:
    "00000000",
    "00000000",
    "00111100",
    "01000010",
    "01111110",
    "01000000",
    "00111100",
    "00000000",


-- # [f] LATIN SMALL LETTER F
-- 0x86:
-- u+0066:
    "00001100",
    "00010010",
    "00010000",
    "01111100",
    "00010000",
    "00010000",
    "00010000",
    "00000000",


-- # [g] LATIN SMALL LETTER G
-- 0x87:
-- u+0067:
    "00000000",
    "00000000",
    "00111010",
    "01000110",
    "01000110",
    "00111010",
    "00000010",
    "00111100",


-- # [h] LATIN SMALL LETTER H
-- 0x88:
-- u+0068:
    "01000000",
    "01000000",
    "01011100",
    "01100010",
    "01000010",
    "01000010",
    "01000010",
    "00000000",


-- # [i] LATIN SMALL LETTER I
-- 0x89:
-- u+0069:
    "00001000",
    "00000000",
    "00011000",
    "00001000",
    "00001000",
    "00001000",
    "00011100",
    "00000000",


-- # [j] LATIN SMALL LETTER J
-- 0x8a:
-- u+006a:
    "00000100",
    "00000000",
    "00001100",
    "00000100",
    "00000100",
    "00000100",
    "01000100",
    "00111000",


-- # [k] LATIN SMALL LETTER K
-- 0x8b:
-- u+006b:
    "01000000",
    "01000000",
    "01000100",
    "01001000",
    "01010000",
    "01101000",
    "01000100",
    "00000000",


-- # [l] LATIN SMALL LETTER L
-- 0x8c:
-- u+006c:
    "00011000",
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00011100",
    "00000000",


-- # [m] LATIN SMALL LETTER M
-- 0x8d:
-- u+006d:
    "00000000",
    "00000000",
    "01110110",
    "01001001",
    "01001001",
    "01001001",
    "01001001",
    "00000000",


-- # [n] LATIN SMALL LETTER N
-- 0x8e:
-- u+006e:
    "00000000",
    "00000000",
    "01011100",
    "01100010",
    "01000010",
    "01000010",
    "01000010",
    "00000000",


-- # [o] LATIN SMALL LETTER O
-- 0x8f:
-- u+006f:
    "00000000",
    "00000000",
    "00111100",
    "01000010",
    "01000010",
    "01000010",
    "00111100",
    "00000000",


-- # [p] LATIN SMALL LETTER P
-- 0x90:
-- u+0070:
    "00000000",
    "00000000",
    "01011100",
    "01100010",
    "01100010",
    "01011100",
    "01000000",
    "01000000",


-- # [q] LATIN SMALL LETTER Q
-- 0x91:
-- u+0071:
    "00000000",
    "00000000",
    "00111010",
    "01000110",
    "01000110",
    "00111010",
    "00000010",
    "00000010",


-- # [r] LATIN SMALL LETTER R
-- 0x92:
-- u+0072:
    "00000000",
    "00000000",
    "01011100",
    "01100010",
    "01000000",
    "01000000",
    "01000000",
    "00000000",


-- # [s] LATIN SMALL LETTER S
-- 0x93:
-- u+0073:
    "00000000",
    "00000000",
    "00111110",
    "01000000",
    "00111100",
    "00000010",
    "01111100",
    "00000000",


-- # [t] LATIN SMALL LETTER T
-- 0x94:
-- u+0074:
    "00010000",
    "00010000",
    "01111100",
    "00010000",
    "00010000",
    "00010010",
    "00001100",
    "00000000",


-- # [u] LATIN SMALL LETTER U
-- 0x95:
-- u+0075:
    "00000000",
    "00000000",
    "01000010",
    "01000010",
    "01000010",
    "01000110",
    "00111010",
    "00000000",


-- # [v] LATIN SMALL LETTER V
-- 0x96:
-- u+0076:
    "00000000",
    "00000000",
    "01000010",
    "01000010",
    "01000010",
    "00100100",
    "00011000",
    "00000000",


-- # [w] LATIN SMALL LETTER W
-- 0x97:
-- u+0077:
    "00000000",
    "00000000",
    "01000001",
    "01001001",
    "01001001",
    "01001001",
    "00110110",
    "00000000",


-- # [x] LATIN SMALL LETTER X
-- 0x98:
-- u+0078:
    "00000000",
    "00000000",
    "01000010",
    "00100100",
    "00011000",
    "00100100",
    "01000010",
    "00000000",


-- # [y] LATIN SMALL LETTER Y
-- 0x99:
-- u+0079:
    "00000000",
    "00000000",
    "01000010",
    "01000010",
    "01000110",
    "00111010",
    "00000010",
    "00111100",


-- # [z] LATIN SMALL LETTER Z
-- 0x9a:
-- u+007a:
    "00000000",
    "00000000",
    "01111110",
    "00000100",
    "00011000",
    "00100000",
    "01111110",
    "00000000",


-- # [[] LEFT SQUARE BRACKET
-- 0x9b:
-- u+005b:
    "00111100",
    "00100000",
    "00100000",
    "00100000",
    "00100000",
    "00100000",
    "00111100",
    "00000000",


-- # [\] REVERSE SOLIDUS
-- 0x9c:
-- u+005c:
    "00000000",
    "01000000",
    "00100000",
    "00010000",
    "00001000",
    "00000100",
    "00000010",
    "00000000",


-- # []] RIGHT SQUARE BRACKET
-- 0x9d:
-- u+005d:
    "00111100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00111100",
    "00000000",


-- # [↑] UPWARDS ARROW
-- 0x9e:
-- u+2191:
    "00000000",
    "00001000",
    "00011100",
    "00101010",
    "00001000",
    "00001000",
    "00001000",
    "00001000",


-- # [←] LEFTWARDS ARROW
-- 0x9f:
-- u+2190:
    "00000000",
    "00000000",
    "00010000",
    "00100000",
    "01111111",
    "00100000",
    "00010000",
    "00000000",


-- # [ ] SPACE
-- 0xa0:
-- u+0020:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",


-- # [!] EXCLAMATION MARK
-- 0xa1:
-- u+0021:
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00000000",
    "00000000",
    "00001000",
    "00000000",


-- # ["] QUOTATION MARK
-- 0xa2:
-- u+0022:
    "00100100",
    "00100100",
    "00100100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",


-- # [-- #] NUMBER SIGN
-- 0xa3:
-- u+0023:
    "00100100",
    "00100100",
    "01111110",
    "00100100",
    "01111110",
    "00100100",
    "00100100",
    "00000000",


-- # [$] DOLLAR SIGN
-- 0xa4:
-- u+0024:
    "00001000",
    "00011110",
    "00101000",
    "00011100",
    "00001010",
    "00111100",
    "00001000",
    "00000000",


-- # [%] PERCENT SIGN
-- 0xa5:
-- u+0025:
    "00000000",
    "01100010",
    "01100100",
    "00001000",
    "00010000",
    "00100110",
    "01000110",
    "00000000",


-- # [&] AMPERSAND
-- 0xa6:
-- u+0026:
    "00110000",
    "01001000",
    "01001000",
    "00110000",
    "01001010",
    "01000100",
    "00111010",
    "00000000",


-- # ['] APOSTROPHE
-- 0xa7:
-- u+0027:
    "00000100",
    "00001000",
    "00010000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",


-- # [(] LEFT PARENTHESIS
-- 0xa8:
-- u+0028:
    "00000100",
    "00001000",
    "00010000",
    "00010000",
    "00010000",
    "00001000",
    "00000100",
    "00000000",


-- # [)] RIGHT PARENTHESIS
-- 0xa9:
-- u+0029:
    "00100000",
    "00010000",
    "00001000",
    "00001000",
    "00001000",
    "00010000",
    "00100000",
    "00000000",


-- # [*] ASTERISK
-- 0xaa:
-- u+002a:
    "00001000",
    "00101010",
    "00011100",
    "00111110",
    "00011100",
    "00101010",
    "00001000",
    "00000000",


-- # [+] PLUS SIGN
-- 0xab:
-- u+002b:
    "00000000",
    "00001000",
    "00001000",
    "00111110",
    "00001000",
    "00001000",
    "00000000",
    "00000000",


-- # [,] COMMA
-- 0xac:
-- u+002c:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00001000",
    "00001000",
    "00010000",


-- # [-] HYPHEN-MINUS
-- 0xad:
-- u+002d:
    "00000000",
    "00000000",
    "00000000",
    "01111110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",


-- # [0] FULL STOP
-- 0xae:
-- u+002e:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011000",
    "00011000",
    "00000000",


-- # [/] SOLIDUS
-- 0xaf:
-- u+002f:
    "00000000",
    "00000010",
    "00000100",
    "00001000",
    "00010000",
    "00100000",
    "01000000",
    "00000000",


-- # [0] DIGIT ZERO
-- 0xb0:
-- u+0030:
    "00111100",
    "01000010",
    "01000110",
    "01011010",
    "01100010",
    "01000010",
    "00111100",
    "00000000",


-- # [1] DIGIT ONE
-- 0xb1:
-- u+0031:
    "00001000",
    "00011000",
    "00101000",
    "00001000",
    "00001000",
    "00001000",
    "00111110",
    "00000000",


-- # [2] DIGIT TWO
-- 0xb2:
-- u+0032:
    "00111100",
    "01000010",
    "00000010",
    "00001100",
    "00110000",
    "01000000",
    "01111110",
    "00000000",


-- # [3] DIGIT THREE
-- 0xb3:
-- u+0033:
    "00111100",
    "01000010",
    "00000010",
    "00011100",
    "00000010",
    "01000010",
    "00111100",
    "00000000",


-- # [4] DIGIT FOUR
-- 0xb4:
-- u+0034:
    "00000100",
    "00001100",
    "00010100",
    "00100100",
    "01111110",
    "00000100",
    "00000100",
    "00000000",


-- # [5] DIGIT FIVE
-- 0xb5:
-- u+0035:
    "01111110",
    "01000000",
    "01111000",
    "00000100",
    "00000010",
    "01000100",
    "00111000",
    "00000000",


-- # [6] DIGIT SIX
-- 0xb6:
-- u+0036:
    "00011100",
    "00100000",
    "01000000",
    "01111100",
    "01000010",
    "01000010",
    "00111100",
    "00000000",


-- # [7] DIGIT SEVEN
-- 0xb7:
-- u+0037:
    "01111110",
    "01000010",
    "00000100",
    "00001000",
    "00010000",
    "00010000",
    "00010000",
    "00000000",


-- # [8] DIGIT EIGHT
-- 0xb8:
-- u+0038:
    "00111100",
    "01000010",
    "01000010",
    "00111100",
    "01000010",
    "01000010",
    "00111100",
    "00000000",


-- # [9] DIGIT NINE
-- 0xb9:
-- u+0039:
    "00111100",
    "01000010",
    "01000010",
    "00111110",
    "00000010",
    "00000100",
    "00111000",
    "00000000",


-- # [:] COLON
-- 0xba:
-- u+003a:
    "00000000",
    "00000000",
    "00001000",
    "00000000",
    "00000000",
    "00001000",
    "00000000",
    "00000000",


-- # [;] SEMICOLON
-- 0xbb:
-- u+003b:
    "00000000",
    "00000000",
    "00001000",
    "00000000",
    "00000000",
    "00001000",
    "00001000",
    "00010000",


-- # [<] LESS-THAN SIGN
-- 0xbc:
-- u+003c:
    "00001110",
    "00011000",
    "00110000",
    "01100000",
    "00110000",
    "00011000",
    "00001110",
    "00000000",


-- # [=] EQUALS SIGN
-- 0xbd:
-- u+003d:
    "00000000",
    "00000000",
    "01111110",
    "00000000",
    "01111110",
    "00000000",
    "00000000",
    "00000000",


-- # [>] GREATER-THAN SIGN
-- 0xbe:
-- u+003e:
    "01110000",
    "00011000",
    "00001100",
    "00000110",
    "00001100",
    "00011000",
    "01110000",
    "00000000",


-- # [?] QUESTION MARK
-- 0xbf:
-- u+003f:
    "00111100",
    "01000010",
    "00000010",
    "00001100",
    "00010000",
    "00000000",
    "00010000",
    "00000000",


-- # [─] BOX DRAWINGS LIGHT HORIZONTAL
-- 0xc0:
-- u+2500:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111111",
    "00000000",
    "00000000",
    "00000000",


-- # [A] LATIN CAPITAL LETTER A
-- 0xc1:
-- u+0041:
    "00011000",
    "00100100",
    "01000010",
    "01111110",
    "01000010",
    "01000010",
    "01000010",
    "00000000",


-- # [B] LATIN CAPITAL LETTER B
-- 0xc2:
-- u+0042:
    "01111100",
    "00100010",
    "00100010",
    "00111100",
    "00100010",
    "00100010",
    "01111100",
    "00000000",


-- # [C] LATIN CAPITAL LETTER C
-- 0xc3:
-- u+0043:
    "00011100",
    "00100010",
    "01000000",
    "01000000",
    "01000000",
    "00100010",
    "00011100",
    "00000000",


-- # [D] LATIN CAPITAL LETTER D
-- 0xc4:
-- u+0044:
    "01111000",
    "00100100",
    "00100010",
    "00100010",
    "00100010",
    "00100100",
    "01111000",
    "00000000",


-- # [E] LATIN CAPITAL LETTER E
-- 0xc5:
-- u+0045:
    "01111110",
    "01000000",
    "01000000",
    "01111000",
    "01000000",
    "01000000",
    "01111110",
    "00000000",


-- # [F] LATIN CAPITAL LETTER F
-- 0xc6:
-- u+0046:
    "01111110",
    "01000000",
    "01000000",
    "01111000",
    "01000000",
    "01000000",
    "01000000",
    "00000000",


-- # [G] LATIN CAPITAL LETTER G
-- 0xc7:
-- u+0047:
    "00011100",
    "00100010",
    "01000000",
    "01001110",
    "01000010",
    "00100010",
    "00011100",
    "00000000",


-- # [H] LATIN CAPITAL LETTER H
-- 0xc8:
-- u+0048:
    "01000010",
    "01000010",
    "01000010",
    "01111110",
    "01000010",
    "01000010",
    "01000010",
    "00000000",


-- # [I] LATIN CAPITAL LETTER I
-- 0xc9:
-- u+0049:
    "00011100",
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00011100",
    "00000000",


-- # [J] LATIN CAPITAL LETTER J
-- 0xca:
-- u+004a:
    "00001110",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "01000100",
    "00111000",
    "00000000",


-- # [K] LATIN CAPITAL LETTER K
-- 0xcb:
-- u+004b:
    "01000010",
    "01000100",
    "01001000",
    "01110000",
    "01001000",
    "01000100",
    "01000010",
    "00000000",


-- # [L] LATIN CAPITAL LETTER L
-- 0xcc:
-- u+004c:
    "01000000",
    "01000000",
    "01000000",
    "01000000",
    "01000000",
    "01000000",
    "01111110",
    "00000000",


-- # [M] LATIN CAPITAL LETTER M
-- 0xcd:
-- u+004d:
    "01000010",
    "01100110",
    "01011010",
    "01011010",
    "01000010",
    "01000010",
    "01000010",
    "00000000",


-- # [N] LATIN CAPITAL LETTER N
-- 0xce:
-- u+004e:
    "01000010",
    "01100010",
    "01010010",
    "01001010",
    "01000110",
    "01000010",
    "01000010",
    "00000000",


-- # [O] LATIN CAPITAL LETTER O
-- 0xcf:
-- u+004f:
    "00011000",
    "00100100",
    "01000010",
    "01000010",
    "01000010",
    "00100100",
    "00011000",
    "00000000",


-- # [P] LATIN CAPITAL LETTER P
-- 0xd0:
-- u+0050:
    "01111100",
    "01000010",
    "01000010",
    "01111100",
    "01000000",
    "01000000",
    "01000000",
    "00000000",


-- # [Q] LATIN CAPITAL LETTER Q
-- 0xd1:
-- u+0051:
    "00011000",
    "00100100",
    "01000010",
    "01000010",
    "01001010",
    "00100100",
    "00011010",
    "00000000",


-- # [R] LATIN CAPITAL LETTER R
-- 0xd2:
-- u+0052:
    "01111100",
    "01000010",
    "01000010",
    "01111100",
    "01001000",
    "01000100",
    "01000010",
    "00000000",


-- # [S] LATIN CAPITAL LETTER S
-- 0xd3:
-- u+0053:
    "00111100",
    "01000010",
    "01000000",
    "00111100",
    "00000010",
    "01000010",
    "00111100",
    "00000000",


-- # [T] LATIN CAPITAL LETTER T
-- 0xd4:
-- u+0054:
    "00111110",
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00000000",


-- # [U] LATIN CAPITAL LETTER U
-- 0xd5:
-- u+0055:
    "01000010",
    "01000010",
    "01000010",
    "01000010",
    "01000010",
    "01000010",
    "00111100",
    "00000000",


-- # [V] LATIN CAPITAL LETTER V
-- 0xd6:
-- u+0056:
    "01000010",
    "01000010",
    "01000010",
    "00100100",
    "00100100",
    "00011000",
    "00011000",
    "00000000",


-- # [W] LATIN CAPITAL LETTER W
-- 0xd7:
-- u+0057:
    "01000010",
    "01000010",
    "01000010",
    "01011010",
    "01011010",
    "01100110",
    "01000010",
    "00000000",


-- # [X] LATIN CAPITAL LETTER X
-- 0xd8:
-- u+0058:
    "01000010",
    "01000010",
    "00100100",
    "00011000",
    "00100100",
    "01000010",
    "01000010",
    "00000000",


-- # [Y] LATIN CAPITAL LETTER Y
-- 0xd9:
-- u+0059:
    "00100010",
    "00100010",
    "00100010",
    "00011100",
    "00001000",
    "00001000",
    "00001000",
    "00000000",


-- # [Z] LATIN CAPITAL LETTER Z
-- 0xda:
-- u+005a:
    "01111110",
    "00000010",
    "00000100",
    "00011000",
    "00100000",
    "01000000",
    "01111110",
    "00000000",


-- # [┼] BOX DRAWINGS LIGHT VERTICAL AND HORIZONTAL
-- 0xdb:
-- u+253c:
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "11111111",
    "00001000",
    "00001000",
    "00001000",


-- # [🮌] LEFT HALF MEDIUM SHADE
-- 0xdc:
-- u+1fb8c:
    "10100000",
    "01010000",
    "10100000",
    "01010000",
    "10100000",
    "01010000",
    "10100000",
    "01010000",


-- # [│] BOX DRAWINGS LIGHT VERTICAL
-- 0xdd:
-- u+2502:
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00001000",


-- # [🮕] CHECKER BOARD FILL
-- 0xde:
-- u+1fb95:
    "11001100",
    "11001100",
    "00110011",
    "00110011",
    "11001100",
    "11001100",
    "00110011",
    "00110011",


-- # [🮘] UPPER LEFT TO LOWER RIGHT FILL
-- 0xdf:
-- u+1fb98:
    "11001100",
    "01100110",
    "00110011",
    "10011001",
    "11001100",
    "01100110",
    "00110011",
    "10011001",


-- # [ ] NO-BREAK SPACE
-- 0xe0:
-- u+00a0:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",


-- # [▌] LEFT HALF BLOCK
-- 0xe1:
-- u+258c:
    "11110000",
    "11110000",
    "11110000",
    "11110000",
    "11110000",
    "11110000",
    "11110000",
    "11110000",


-- # [▄] LOWER HALF BLOCK
-- 0xe2:
-- u+2584:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111111",
    "11111111",
    "11111111",
    "11111111",


-- # [▔] UPPER ONE EIGHTH BLOCK
-- 0xe3:
-- u+2594:
    "11111111",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",


-- # [▁] LOWER ONE EIGHTH BLOCK
-- 0xe4:
-- u+2581:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111111",


-- # [▏] LEFT ONE EIGHTH BLOCK
-- 0xe5:
-- u+258f:
    "10000000",
    "10000000",
    "10000000",
    "10000000",
    "10000000",
    "10000000",
    "10000000",
    "10000000",


-- # [▒] MEDIUM SHADE
-- 0xe6:
-- u+2592:
    "10101010",
    "01010101",
    "10101010",
    "01010101",
    "10101010",
    "01010101",
    "10101010",
    "01010101",


-- # [▕] RIGHT ONE EIGHTH BLOCK
-- 0xe7:
-- u+2595:
    "00000001",
    "00000001",
    "00000001",
    "00000001",
    "00000001",
    "00000001",
    "00000001",
    "00000001",


-- # [🮏] LOWER HALF MEDIUM SHADE
-- 0xe8:
-- u+1fb8f:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "10101010",
    "01010101",
    "10101010",
    "01010101",


-- # [🮙] UPPER RIGHT TO LOWER LEFT FILL
-- 0xe9:
-- u+1fb99:
    "10011001",
    "00110011",
    "01100110",
    "11001100",
    "10011001",
    "00110011",
    "01100110",
    "11001100",


-- # [🮇] RIGHT ONE QUARTER BLOCK
-- 0xea:
-- u+1fb87:
    "00000011",
    "00000011",
    "00000011",
    "00000011",
    "00000011",
    "00000011",
    "00000011",
    "00000011",


-- # [├] BOX DRAWINGS LIGHT VERTICAL AND RIGHT
-- 0xeb:
-- u+251c:
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00001111",
    "00001000",
    "00001000",
    "00001000",


-- # [▗] QUADRANT LOWER RIGHT
-- 0xec:
-- u+2597:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00001111",
    "00001111",
    "00001111",
    "00001111",


-- # [└] BOX DRAWINGS LIGHT UP AND RIGHT
-- 0xed:
-- u+2514:
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00001111",
    "00000000",
    "00000000",
    "00000000",


-- # [┐] BOX DRAWINGS LIGHT DOWN AND LEFT
-- 0xee:
-- u+2510:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111000",
    "00001000",
    "00001000",
    "00001000",


-- # [▂] LOWER ONE QUARTER BLOCK
-- 0xef:
-- u+2582:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111111",
    "11111111",


-- # [┌] BOX DRAWINGS LIGHT DOWN AND RIGHT
-- 0xf0:
-- u+250c:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00001111",
    "00001000",
    "00001000",
    "00001000",


-- # [┴] BOX DRAWINGS LIGHT UP AND HORIZONTAL
-- 0xf1:
-- u+2534:
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "11111111",
    "00000000",
    "00000000",
    "00000000",


-- # [┬] BOX DRAWINGS LIGHT DOWN AND HORIZONTAL
-- 0xf2:
-- u+252c:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111111",
    "00001000",
    "00001000",
    "00001000",


-- # [┤] BOX DRAWINGS LIGHT VERTICAL AND LEFT
-- 0xf3:
-- u+2524:
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "11111000",
    "00001000",
    "00001000",
    "00001000",


-- # [▎] LEFT ONE QUARTER BLOCK
-- 0xf4:
-- u+258e:
    "11000000",
    "11000000",
    "11000000",
    "11000000",
    "11000000",
    "11000000",
    "11000000",
    "11000000",


-- # [▍] LEFT THREE EIGHTHS BLOCK
-- 0xf5:
-- u+258d:
    "11100000",
    "11100000",
    "11100000",
    "11100000",
    "11100000",
    "11100000",
    "11100000",
    "11100000",


-- # [🮈] RIGHT THREE EIGHTHS BLOCK
-- 0xf6:
-- u+1fb88:
    "00000111",
    "00000111",
    "00000111",
    "00000111",
    "00000111",
    "00000111",
    "00000111",
    "00000111",


-- # [🮂] UPPER ONE QUARTER BLOCK
-- 0xf7:
-- u+1fb82:
    "11111111",
    "11111111",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",


-- # [🮃] UPPER THREE EIGHTHS BLOCK
-- 0xf8:
-- u+1fb83:
    "11111111",
    "11111111",
    "11111111",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",


-- # [▃] LOWER THREE EIGHTHS BLOCK
-- 0xf9:
-- u+2583:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111111",
    "11111111",
    "11111111",


-- # [✓] CHECK MARK
-- 0xfa:
-- u+2713:
    "00000001",
    "00000010",
    "01000100",
    "01001000",
    "01010000",
    "01100000",
    "01000000",
    "00000000",


-- # [▖] QUADRANT LOWER LEFT
-- 0xfb:
-- u+2596:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11110000",
    "11110000",
    "11110000",
    "11110000",


-- # [▝] QUADRANT UPPER RIGHT
-- 0xfc:
-- u+259d:
    "00001111",
    "00001111",
    "00001111",
    "00001111",
    "00000000",
    "00000000",
    "00000000",
    "00000000",


-- # [┘] BOX DRAWINGS LIGHT UP AND LEFT
-- 0xfd:
-- u+2518:
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "11111000",
    "00000000",
    "00000000",
    "00000000",


-- # [▘] QUADRANT UPPER LEFT
-- 0xfe:
-- u+2598:
    "11110000",
    "11110000",
    "11110000",
    "11110000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",


-- # [▚] QUADRANT UPPER LEFT AND LOWER RIGHT
-- 0xff:
-- u+259a:
    "11110000",
    "11110000",
    "11110000",
    "11110000",
    "00001111",
    "00001111",
    "00001111",
    "00001111",

    );
begin

    dataOut <= ROM(to_integer(unsigned(addrIn)));

end architecture rtl;