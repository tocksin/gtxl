-- @file rom_font.vhd
-- @brief ROM containing character font
-- @author Justin Davis
--
-- $Revision: -
-- $Date: 06/22/2023
-- $LastEditedBy: Justin Davis
--
-- Developed by 2023 Southwest Research Institute
-------------------------------------------------------------------------------
-- Font data taken from: https://github.com/robhagemans/hoard-of-bitfonts/blob/master/commodore/pet/pet.yaff

library ieee;           use ieee.std_logic_1164.all;
                        use ieee.numeric_std.all;

library work;           use work.tools_pkg.all;
                        use work.sys_description_pkg.all;

entity rom_font is
    port ( addrIn   : in    slv(10 downto 0) ;
           dataOut  :   out slv(7 downto 0));
end entity rom_font;

architecture rtl of rom_font is
   
    type rom_type is array (0 to (2**addrIn'length)-1) of std_logic_vector(dataOut'range);

    -- ROM definition
    signal rom : rom_type := ( 

-- 0x00:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00111110",
    "00111110",
    "00111110",
    "00111110",

-- 0x01:
-- u+2502:
    "00010000",
    "00010000",
    "00010000",
    "00010000",
    "00010000",
    "00010000",
    "00010000",
    "00010000",

-- 0x02:
-- u+2500:
    "00000000",
    "00000000",
    "00000000",
    "11111111",
    "00000000",
    "00000000",
    "00000000",
    "00000000",

-- 0x03:
-- u+2518:
    "00010000",
    "00010000",
    "00010000",
    "11110000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",

-- 0x04:
-- u+2514:
    "00010000",
    "00010000",
    "00010000",
    "00011111",
    "00000000",
    "00000000",
    "00000000",
    "00000000",

-- 0x05:
-- u+250c:
    "00000000",
    "00000000",
    "00000000",
    "00011111",
    "00010000",
    "00010000",
    "00010000",
    "00010000",

-- 0x06:
-- u+2510:
    "00000000",
    "00000000",
    "00000000",
    "11110000",
    "00010000",
    "00010000",
    "00010000",
    "00010000",

-- 0x07:
-- u+2534:
    "00010000",
    "00010000",
    "00010000",
    "11111111",
    "00000000",
    "00000000",
    "00000000",
    "00000000",

-- 0x08:
-- u+251c:
    "00010000",
    "00010000",
    "00010000",
    "00011111",
    "00010000",
    "00010000",
    "00010000",
    "00010000",

-- 0x09:
-- u+252c:
    "00000000",
    "00000000",
    "00000000",
    "11111111",
    "00010000",
    "00010000",
    "00010000",
    "00010000",

-- 0x0a:
-- u+2524:
    "00010000",
    "00010000",
    "00010000",
    "11110000",
    "00010000",
    "00010000",
    "00010000",
    "00010000",

-- 0x0b:
-- u+253c:
    "00010000",
    "00010000",
    "00010000",
    "11111111",
    "00010000",
    "00010000",
    "00010000",
    "00010000",

-- 0x0c:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00111110",
    "00111110",
    "00111110",
    "00111110",

-- 0x0d:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00111110",
    "00111110",
    "00111110",
    "00111110",

-- 0x0e:
-- u+2371:
    "00100000",
    "01010100",
    "00001000",
    "00000000",
    "01000100",
    "00101000",
    "00010000",
    "00000000",

-- 0x0f:
-- u+2372:
    "00100000",
    "01010100",
    "00001000",
    "00000000",
    "00010000",
    "00101000",
    "01000100",
    "00000000",

-- 0x10:
-- u+2352:
    "00010000",
    "00010000",
    "01111100",
    "01010100",
    "00101000",
    "00010000",
    "00010000",
    "00000000",

-- 0x11:
-- u+234b:
    "00010000",
    "00010000",
    "00101000",
    "01010100",
    "01111100",
    "00010000",
    "00010000",
    "00000000",

-- 0x12:
-- u+233d:
    "00010000",
    "00111000",
    "01010100",
    "01010100",
    "01010100",
    "00111000",
    "00010000",
    "00000000",

-- 0x13:
-- u+2349:
    "10000000",
    "01111000",
    "01100100",
    "01010100",
    "01001100",
    "00111100",
    "00000010",
    "00000000",

-- 0x14:
-- u+2296:
    "00000000",
    "00111000",
    "01000100",
    "11111110",
    "01000100",
    "00111000",
    "00000000",
    "00000000",

-- 0x15:
-- u+2295:
    "00000000",
    "00111000",
    "01010100",
    "01111100",
    "01010100",
    "00111000",
    "00000000",
    "00000000",

-- 0x16:
-- u+236b:
    "00100000",
    "01010100",
    "00001000",
    "00000000",
    "01111100",
    "01000100",
    "00101000",
    "00010000",

-- 0x17:
-- u+234e:
    "00000000",
    "00000000",
    "00111000",
    "00101000",
    "00111000",
    "00010000",
    "01111100",
    "00000000",

-- 0x18:
-- u+2355:
    "00000000",
    "00000000",
    "01111100",
    "00010000",
    "00111000",
    "00101000",
    "00111000",
    "00000000",

-- 0x19:
-- u+2340:
    "00000000",
    "01000000",
    "00100000",
    "01111100",
    "00001000",
    "00000100",
    "00000010",
    "00000000",

-- 0x1a:
-- u+233f:
    "00000000",
    "00000100",
    "00001000",
    "01111100",
    "00100000",
    "01000000",
    "10000000",
    "00000000",

-- 0x1b:
-- u+235d:
    "00000000",
    "00000000",
    "00110000",
    "01001000",
    "01001000",
    "01111000",
    "01001000",
    "00000000",

-- 0x1c:
-- u+235e:
    "01111100",
    "01010100",
    "01010100",
    "01000100",
    "01000100",
    "01000100",
    "01111100",
    "00000000",

-- 0x1d:
-- u+0021:
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00000000",
    "00000000",
    "00001000",
    "00000000",

-- 0x1e:
-- u+2339:
    "01111100",
    "01010100",
    "01000100",
    "01111100",
    "01000100",
    "01010100",
    "01111100",
    "00000000",

-- 0x1f:
-- u+2336:
    "00000000",
    "00000000",
    "01111100",
    "00010000",
    "00010000",
    "00010000",
    "01111100",
    "00000000",

-- # [ ] SPACE
-- 0x20:
-- u+0020:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",


-- # [!] EXCLAMATION MARK
-- 0x21:
-- u+0021:
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00000000",
    "00000000",
    "00001000",
    "00000000",


-- # ["] QUOTATION MARK
-- 0x22:
-- u+0022:
    "00100100",
    "00100100",
    "00100100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",


-- # [-- #] NUMBER SIGN
-- 0x23:
-- u+0023:
    "00100100",
    "00100100",
    "01111110",
    "00100100",
    "01111110",
    "00100100",
    "00100100",
    "00000000",


-- # [$] DOLLAR SIGN
-- 0x24:
-- u+0024:
    "00001000",
    "00011110",
    "00101000",
    "00011100",
    "00001010",
    "00111100",
    "00001000",
    "00000000",


-- # [%] PERCENT SIGN
-- 0x25:
-- u+0025:
    "00000000",
    "01100010",
    "01100100",
    "00001000",
    "00010000",
    "00100110",
    "01000110",
    "00000000",


-- # [&] AMPERSAND
-- 0x26:
-- u+0026:
    "00110000",
    "01001000",
    "01001000",
    "00110000",
    "01001010",
    "01000100",
    "00111010",
    "00000000",


-- # ['] APOSTROPHE
-- 0x27:
-- u+0027:
    "00000100",
    "00001000",
    "00010000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",


-- # [(] LEFT PARENTHESIS
-- 0x28:
-- u+0028:
    "00000100",
    "00001000",
    "00010000",
    "00010000",
    "00010000",
    "00001000",
    "00000100",
    "00000000",


-- # [)] RIGHT PARENTHESIS
-- 0x29:
-- u+0029:
    "00100000",
    "00010000",
    "00001000",
    "00001000",
    "00001000",
    "00010000",
    "00100000",
    "00000000",


-- # [*] ASTERISK
-- 0x2a:
-- u+002a:
    "00001000",
    "00101010",
    "00011100",
    "00111110",
    "00011100",
    "00101010",
    "00001000",
    "00000000",


-- # [+] PLUS SIGN
-- 0x2b:
-- u+002b:
    "00000000",
    "00001000",
    "00001000",
    "00111110",
    "00001000",
    "00001000",
    "00000000",
    "00000000",


-- # [,] COMMA
-- 0x2c:
-- u+002c:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00001000",
    "00001000",
    "00010000",


-- # [-] HYPHEN-MINUS
-- 0x2d:
-- u+002d:
    "00000000",
    "00000000",
    "00000000",
    "01111110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",


-- # [0] FULL STOP
-- 0x2e:
-- u+002e:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011000",
    "00011000",
    "00000000",


-- # [/] SOLIDUS
-- 0x2f:
-- u+002f:
    "00000000",
    "00000010",
    "00000100",
    "00001000",
    "00010000",
    "00100000",
    "01000000",
    "00000000",


-- # [0] DIGIT ZERO
-- 0x30:
-- u+0030:
    "00111100",
    "01000010",
    "01000110",
    "01011010",
    "01100010",
    "01000010",
    "00111100",
    "00000000",


-- # [1] DIGIT ONE
-- 0x31:
-- u+0031:
    "00001000",
    "00011000",
    "00101000",
    "00001000",
    "00001000",
    "00001000",
    "00111110",
    "00000000",


-- # [2] DIGIT TWO
-- 0x32:
-- u+0032:
    "00111100",
    "01000010",
    "00000010",
    "00001100",
    "00110000",
    "01000000",
    "01111110",
    "00000000",


-- # [3] DIGIT THREE
-- 0x33:
-- u+0033:
    "00111100",
    "01000010",
    "00000010",
    "00011100",
    "00000010",
    "01000010",
    "00111100",
    "00000000",


-- # [4] DIGIT FOUR
-- 0x34:
-- u+0034:
    "00000100",
    "00001100",
    "00010100",
    "00100100",
    "01111110",
    "00000100",
    "00000100",
    "00000000",


-- # [5] DIGIT FIVE
-- 0x35:
-- u+0035:
    "01111110",
    "01000000",
    "01111000",
    "00000100",
    "00000010",
    "01000100",
    "00111000",
    "00000000",


-- # [6] DIGIT SIX
-- 0x36:
-- u+0036:
    "00011100",
    "00100000",
    "01000000",
    "01111100",
    "01000010",
    "01000010",
    "00111100",
    "00000000",


-- # [7] DIGIT SEVEN
-- 0x37:
-- u+0037:
    "01111110",
    "01000010",
    "00000100",
    "00001000",
    "00010000",
    "00010000",
    "00010000",
    "00000000",


-- # [8] DIGIT EIGHT
-- 0x38:
-- u+0038:
    "00111100",
    "01000010",
    "01000010",
    "00111100",
    "01000010",
    "01000010",
    "00111100",
    "00000000",


-- # [9] DIGIT NINE
-- 0x39:
-- u+0039:
    "00111100",
    "01000010",
    "01000010",
    "00111110",
    "00000010",
    "00000100",
    "00111000",
    "00000000",


-- # [:] COLON
-- 0x3a:
-- u+003a:
    "00000000",
    "00000000",
    "00001000",
    "00000000",
    "00000000",
    "00001000",
    "00000000",
    "00000000",


-- # [;] SEMICOLON
-- 0x3b:
-- u+003b:
    "00000000",
    "00000000",
    "00001000",
    "00000000",
    "00000000",
    "00001000",
    "00001000",
    "00010000",


-- # [<] LESS-THAN SIGN
-- 0x3c:
-- u+003c:
    "00001110",
    "00011000",
    "00110000",
    "01100000",
    "00110000",
    "00011000",
    "00001110",
    "00000000",


-- # [=] EQUALS SIGN
-- 0x3d:
-- u+003d:
    "00000000",
    "00000000",
    "01111110",
    "00000000",
    "01111110",
    "00000000",
    "00000000",
    "00000000",


-- # [>] GREATER-THAN SIGN
-- 0x3e:
-- u+003e:
    "01110000",
    "00011000",
    "00001100",
    "00000110",
    "00001100",
    "00011000",
    "01110000",
    "00000000",


-- # [?] QUESTION MARK
-- 0x3f:
-- u+003f:
    "00111100",
    "01000010",
    "00000010",
    "00001100",
    "00010000",
    "00000000",
    "00010000",
    "00000000",


-- # [1] COMMERCIAL AT
-- 0x40:
-- u+0040:
    "00011100",
    "00100010",
    "01001010",
    "01010110",
    "01001100",
    "00100000",
    "00011110",
    "00000000",


-- # [A] LATIN CAPITAL LETTER A
-- 0x41:
-- u+0041:
    "00011000",
    "00100100",
    "01000010",
    "01111110",
    "01000010",
    "01000010",
    "01000010",
    "00000000",


-- # [B] LATIN CAPITAL LETTER B
-- 0x42:
-- u+0042:
    "01111100",
    "00100010",
    "00100010",
    "00111100",
    "00100010",
    "00100010",
    "01111100",
    "00000000",


-- # [C] LATIN CAPITAL LETTER C
-- 0x43:
-- u+0043:
    "00011100",
    "00100010",
    "01000000",
    "01000000",
    "01000000",
    "00100010",
    "00011100",
    "00000000",


-- # [D] LATIN CAPITAL LETTER D
-- 0x44:
-- u+0044:
    "01111000",
    "00100100",
    "00100010",
    "00100010",
    "00100010",
    "00100100",
    "01111000",
    "00000000",


-- # [E] LATIN CAPITAL LETTER E
-- 0x45:
-- u+0045:
    "01111110",
    "01000000",
    "01000000",
    "01111000",
    "01000000",
    "01000000",
    "01111110",
    "00000000",


-- # [F] LATIN CAPITAL LETTER F
-- 0x46:
-- u+0046:
    "01111110",
    "01000000",
    "01000000",
    "01111000",
    "01000000",
    "01000000",
    "01000000",
    "00000000",


-- # [G] LATIN CAPITAL LETTER G
-- 0x47:
-- u+0047:
    "00011100",
    "00100010",
    "01000000",
    "01001110",
    "01000010",
    "00100010",
    "00011100",
    "00000000",


-- # [H] LATIN CAPITAL LETTER H
-- 0x48:
-- u+0048:
    "01000010",
    "01000010",
    "01000010",
    "01111110",
    "01000010",
    "01000010",
    "01000010",
    "00000000",


-- # [I] LATIN CAPITAL LETTER I
-- 0x49:
-- u+0049:
    "00011100",
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00011100",
    "00000000",


-- # [J] LATIN CAPITAL LETTER J
-- 0x4a:
-- u+004a:
    "00001110",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "01000100",
    "00111000",
    "00000000",


-- # [K] LATIN CAPITAL LETTER K
-- 0x4b:
-- u+004b:
    "01000010",
    "01000100",
    "01001000",
    "01110000",
    "01001000",
    "01000100",
    "01000010",
    "00000000",


-- # [L] LATIN CAPITAL LETTER L
-- 0x4c:
-- u+004c:
    "01000000",
    "01000000",
    "01000000",
    "01000000",
    "01000000",
    "01000000",
    "01111110",
    "00000000",


-- # [M] LATIN CAPITAL LETTER M
-- 0x4d:
-- u+004d:
    "01000010",
    "01100110",
    "01011010",
    "01011010",
    "01000010",
    "01000010",
    "01000010",
    "00000000",


-- # [N] LATIN CAPITAL LETTER N
-- 0x4e:
-- u+004e:
    "01000010",
    "01100010",
    "01010010",
    "01001010",
    "01000110",
    "01000010",
    "01000010",
    "00000000",


-- # [O] LATIN CAPITAL LETTER O
-- 0x4f:
-- u+004f:
    "00011000",
    "00100100",
    "01000010",
    "01000010",
    "01000010",
    "00100100",
    "00011000",
    "00000000",


-- # [P] LATIN CAPITAL LETTER P
-- 0x50:
-- u+0050:
    "01111100",
    "01000010",
    "01000010",
    "01111100",
    "01000000",
    "01000000",
    "01000000",
    "00000000",


-- # [Q] LATIN CAPITAL LETTER Q
-- 0x51:
-- u+0051:
    "00011000",
    "00100100",
    "01000010",
    "01000010",
    "01001010",
    "00100100",
    "00011010",
    "00000000",


-- # [R] LATIN CAPITAL LETTER R
-- 0x52:
-- u+0052:
    "01111100",
    "01000010",
    "01000010",
    "01111100",
    "01001000",
    "01000100",
    "01000010",
    "00000000",


-- # [S] LATIN CAPITAL LETTER S
-- 0x53:
-- u+0053:
    "00111100",
    "01000010",
    "01000000",
    "00111100",
    "00000010",
    "01000010",
    "00111100",
    "00000000",


-- # [T] LATIN CAPITAL LETTER T
-- 0x54:
-- u+0054:
    "00111110",
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00000000",


-- # [U] LATIN CAPITAL LETTER U
-- 0x55:
-- u+0055:
    "01000010",
    "01000010",
    "01000010",
    "01000010",
    "01000010",
    "01000010",
    "00111100",
    "00000000",


-- # [V] LATIN CAPITAL LETTER V
-- 0x56:
-- u+0056:
    "01000010",
    "01000010",
    "01000010",
    "00100100",
    "00100100",
    "00011000",
    "00011000",
    "00000000",


-- # [W] LATIN CAPITAL LETTER W
-- 0x57:
-- u+0057:
    "01000010",
    "01000010",
    "01000010",
    "01011010",
    "01011010",
    "01100110",
    "01000010",
    "00000000",


-- # [X] LATIN CAPITAL LETTER X
-- 0x58:
-- u+0058:
    "01000010",
    "01000010",
    "00100100",
    "00011000",
    "00100100",
    "01000010",
    "01000010",
    "00000000",


-- # [Y] LATIN CAPITAL LETTER Y
-- 0x59:
-- u+0059:
    "00100010",
    "00100010",
    "00100010",
    "00011100",
    "00001000",
    "00001000",
    "00001000",
    "00000000",


-- # [Z] LATIN CAPITAL LETTER Z
-- 0x5a:
-- u+005a:
    "01111110",
    "00000010",
    "00000100",
    "00011000",
    "00100000",
    "01000000",
    "01111110",
    "00000000",


-- # [[] LEFT SQUARE BRACKET
-- 0x5b:
-- u+005b:
    "00111100",
    "00100000",
    "00100000",
    "00100000",
    "00100000",
    "00100000",
    "00111100",
    "00000000",


-- # [\] REVERSE SOLIDUS
-- 0x5c:
-- u+005c:
    "00000000",
    "01000000",
    "00100000",
    "00010000",
    "00001000",
    "00000100",
    "00000010",
    "00000000",


-- # []] RIGHT SQUARE BRACKET
-- 0x5d:
-- u+005d:
    "00111100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00111100",
    "00000000",


-- # [^] CIRCUMFLEX ACCENT
-- 0x5e:
-- u+005e:
    "00010000",
    "00101000",
    "01000100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",


-- # [_] LOW LINE
-- 0x5f:
-- u+005f:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111110",


-- # [`] GRAVE ACCENT
-- 0x60:
-- u+0060:
    "00100000",
    "00010000",
    "00001000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",


-- # [a] LATIN SMALL LETTER A
-- 0x61:
-- u+0061:
    "00000000",
    "00000000",
    "00111000",
    "00000100",
    "00111100",
    "01000100",
    "00111010",
    "00000000",


-- # [b] LATIN SMALL LETTER B
-- 0x62:
-- u+0062:
    "01000000",
    "01000000",
    "01011100",
    "01100010",
    "01000010",
    "01100010",
    "01011100",
    "00000000",


-- # [c] LATIN SMALL LETTER C
-- 0x63:
-- u+0063:
    "00000000",
    "00000000",
    "00111100",
    "01000010",
    "01000000",
    "01000010",
    "00111100",
    "00000000",


-- # [d] LATIN SMALL LETTER D
-- 0x64:
-- u+0064:
    "00000010",
    "00000010",
    "00111010",
    "01000110",
    "01000010",
    "01000110",
    "00111010",
    "00000000",


-- # [e] LATIN SMALL LETTER E
-- 0x65:
-- u+0065:
    "00000000",
    "00000000",
    "00111100",
    "01000010",
    "01111110",
    "01000000",
    "00111100",
    "00000000",


-- # [f] LATIN SMALL LETTER F
-- 0x66:
-- u+0066:
    "00001100",
    "00010010",
    "00010000",
    "01111100",
    "00010000",
    "00010000",
    "00010000",
    "00000000",


-- # [g] LATIN SMALL LETTER G
-- 0x67:
-- u+0067:
    "00000000",
    "00000000",
    "00111010",
    "01000110",
    "01000110",
    "00111010",
    "00000010",
    "00111100",


-- # [h] LATIN SMALL LETTER H
-- 0x68:
-- u+0068:
    "01000000",
    "01000000",
    "01011100",
    "01100010",
    "01000010",
    "01000010",
    "01000010",
    "00000000",


-- # [i] LATIN SMALL LETTER I
-- 0x69:
-- u+0069:
    "00001000",
    "00000000",
    "00011000",
    "00001000",
    "00001000",
    "00001000",
    "00011100",
    "00000000",


-- # [j] LATIN SMALL LETTER J
-- 0x6a:
-- u+006a:
    "00000100",
    "00000000",
    "00001100",
    "00000100",
    "00000100",
    "00000100",
    "01000100",
    "00111000",


-- # [k] LATIN SMALL LETTER K
-- 0x6b:
-- u+006b:
    "01000000",
    "01000000",
    "01000100",
    "01001000",
    "01010000",
    "01101000",
    "01000100",
    "00000000",


-- # [l] LATIN SMALL LETTER L
-- 0x6c:
-- u+006c:
    "00011000",
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00011100",
    "00000000",


-- # [m] LATIN SMALL LETTER M
-- 0x6d:
-- u+006d:
    "00000000",
    "00000000",
    "01110110",
    "01001001",
    "01001001",
    "01001001",
    "01001001",
    "00000000",


-- # [n] LATIN SMALL LETTER N
-- 0x6e:
-- u+006e:
    "00000000",
    "00000000",
    "01011100",
    "01100010",
    "01000010",
    "01000010",
    "01000010",
    "00000000",


-- # [o] LATIN SMALL LETTER O
-- 0x6f:
-- u+006f:
    "00000000",
    "00000000",
    "00111100",
    "01000010",
    "01000010",
    "01000010",
    "00111100",
    "00000000",


-- # [p] LATIN SMALL LETTER P
-- 0x70:
-- u+0070:
    "00000000",
    "00000000",
    "01011100",
    "01100010",
    "01100010",
    "01011100",
    "01000000",
    "01000000",


-- # [q] LATIN SMALL LETTER Q
-- 0x71:
-- u+0071:
    "00000000",
    "00000000",
    "00111010",
    "01000110",
    "01000110",
    "00111010",
    "00000010",
    "00000010",


-- # [r] LATIN SMALL LETTER R
-- 0x72:
-- u+0072:
    "00000000",
    "00000000",
    "01011100",
    "01100010",
    "01000000",
    "01000000",
    "01000000",
    "00000000",


-- # [s] LATIN SMALL LETTER S
-- 0x73:
-- u+0073:
    "00000000",
    "00000000",
    "00111110",
    "01000000",
    "00111100",
    "00000010",
    "01111100",
    "00000000",


-- # [t] LATIN SMALL LETTER T
-- 0x74:
-- u+0074:
    "00010000",
    "00010000",
    "01111100",
    "00010000",
    "00010000",
    "00010010",
    "00001100",
    "00000000",


-- # [u] LATIN SMALL LETTER U
-- 0x75:
-- u+0075:
    "00000000",
    "00000000",
    "01000010",
    "01000010",
    "01000010",
    "01000110",
    "00111010",
    "00000000",


-- # [v] LATIN SMALL LETTER V
-- 0x76:
-- u+0076:
    "00000000",
    "00000000",
    "01000010",
    "01000010",
    "01000010",
    "00100100",
    "00011000",
    "00000000",


-- # [w] LATIN SMALL LETTER W
-- 0x77:
-- u+0077:
    "00000000",
    "00000000",
    "01000001",
    "01001001",
    "01001001",
    "01001001",
    "00110110",
    "00000000",


-- # [x] LATIN SMALL LETTER X
-- 0x78:
-- u+0078:
    "00000000",
    "00000000",
    "01000010",
    "00100100",
    "00011000",
    "00100100",
    "01000010",
    "00000000",


-- # [y] LATIN SMALL LETTER Y
-- 0x79:
-- u+0079:
    "00000000",
    "00000000",
    "01000010",
    "01000010",
    "01000110",
    "00111010",
    "00000010",
    "00111100",


-- # [z] LATIN SMALL LETTER Z
-- 0x7a:
-- u+007a:
    "00000000",
    "00000000",
    "01111110",
    "00000100",
    "00011000",
    "00100000",
    "01111110",
    "00000000",


-- # [{] LEFT CURLY BRACKET
-- 0x7b:
-- u+007b:
    "00011000",
    "00100000",
    "00100000",
    "01000000",
    "00100000",
    "00100000",
    "00011000",
    "00000000",


-- # [|] VERTICAL LINE
-- 0x7c:
-- u+007c:
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00001000",


-- # [}] RIGHT CURLY BRACKET
-- 0x7d:
-- u+007d:
    "00110000",
    "00001000",
    "00001000",
    "00000100",
    "00001000",
    "00001000",
    "00110000",
    "00000000",


-- # [~] TILDE
-- 0x7e:
-- u+007e:
    "00000000",
    "00000000",
    "00000000",
    "00100000",
    "01010100",
    "00001000",
    "00000000",
    "00000000",

-- 0x7f:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00111110",
    "00111110",
    "00111110",
    "00111110",

-- 0x00:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00111110",
    "00111110",
    "00111110",
    "00111110",

-- 0x01:
-- u+2502:
    "00010000",
    "00010000",
    "00010000",
    "00010000",
    "00010000",
    "00010000",
    "00010000",
    "00010000",

-- 0x02:
-- u+2500:
    "00000000",
    "00000000",
    "00000000",
    "11111111",
    "00000000",
    "00000000",
    "00000000",
    "00000000",

-- 0x03:
-- u+2518:
    "00010000",
    "00010000",
    "00010000",
    "11110000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",

-- 0x04:
-- u+2514:
    "00010000",
    "00010000",
    "00010000",
    "00011111",
    "00000000",
    "00000000",
    "00000000",
    "00000000",

-- 0x05:
-- u+250c:
    "00000000",
    "00000000",
    "00000000",
    "00011111",
    "00010000",
    "00010000",
    "00010000",
    "00010000",

-- 0x06:
-- u+2510:
    "00000000",
    "00000000",
    "00000000",
    "11110000",
    "00010000",
    "00010000",
    "00010000",
    "00010000",

-- 0x07:
-- u+2534:
    "00010000",
    "00010000",
    "00010000",
    "11111111",
    "00000000",
    "00000000",
    "00000000",
    "00000000",

-- 0x08:
-- u+251c:
    "00010000",
    "00010000",
    "00010000",
    "00011111",
    "00010000",
    "00010000",
    "00010000",
    "00010000",

-- 0x09:
-- u+252c:
    "00000000",
    "00000000",
    "00000000",
    "11111111",
    "00010000",
    "00010000",
    "00010000",
    "00010000",

-- 0x0a:
-- u+2524:
    "00010000",
    "00010000",
    "00010000",
    "11110000",
    "00010000",
    "00010000",
    "00010000",
    "00010000",

-- 0x0b:
-- u+253c:
    "00010000",
    "00010000",
    "00010000",
    "11111111",
    "00010000",
    "00010000",
    "00010000",
    "00010000",

-- 0x0c:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00111110",
    "00111110",
    "00111110",
    "00111110",

-- 0x0d:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00111110",
    "00111110",
    "00111110",
    "00111110",

-- 0x0e:
-- u+2371:
    "00100000",
    "01010100",
    "00001000",
    "00000000",
    "01000100",
    "00101000",
    "00010000",
    "00000000",

-- 0x0f:
-- u+2372:
    "00100000",
    "01010100",
    "00001000",
    "00000000",
    "00010000",
    "00101000",
    "01000100",
    "00000000",

-- 0x10:
-- u+2352:
    "00010000",
    "00010000",
    "01111100",
    "01010100",
    "00101000",
    "00010000",
    "00010000",
    "00000000",

-- 0x11:
-- u+234b:
    "00010000",
    "00010000",
    "00101000",
    "01010100",
    "01111100",
    "00010000",
    "00010000",
    "00000000",

-- 0x12:
-- u+233d:
    "00010000",
    "00111000",
    "01010100",
    "01010100",
    "01010100",
    "00111000",
    "00010000",
    "00000000",

-- 0x13:
-- u+2349:
    "10000000",
    "01111000",
    "01100100",
    "01010100",
    "01001100",
    "00111100",
    "00000010",
    "00000000",

-- 0x14:
-- u+2296:
    "00000000",
    "00111000",
    "01000100",
    "11111110",
    "01000100",
    "00111000",
    "00000000",
    "00000000",

-- 0x15:
-- u+2295:
    "00000000",
    "00111000",
    "01010100",
    "01111100",
    "01010100",
    "00111000",
    "00000000",
    "00000000",

-- 0x16:
-- u+236b:
    "00100000",
    "01010100",
    "00001000",
    "00000000",
    "01111100",
    "01000100",
    "00101000",
    "00010000",

-- 0x17:
-- u+234e:
    "00000000",
    "00000000",
    "00111000",
    "00101000",
    "00111000",
    "00010000",
    "01111100",
    "00000000",

-- 0x18:
-- u+2355:
    "00000000",
    "00000000",
    "01111100",
    "00010000",
    "00111000",
    "00101000",
    "00111000",
    "00000000",

-- 0x19:
-- u+2340:
    "00000000",
    "01000000",
    "00100000",
    "01111100",
    "00001000",
    "00000100",
    "00000010",
    "00000000",

-- 0x1a:
-- u+233f:
    "00000000",
    "00000100",
    "00001000",
    "01111100",
    "00100000",
    "01000000",
    "10000000",
    "00000000",

-- 0x1b:
-- u+235d:
    "00000000",
    "00000000",
    "00110000",
    "01001000",
    "01001000",
    "01111000",
    "01001000",
    "00000000",

-- 0x1c:
-- u+235e:
    "01111100",
    "01010100",
    "01010100",
    "01000100",
    "01000100",
    "01000100",
    "01111100",
    "00000000",

-- 0x1d:
-- u+0021:
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00000000",
    "00000000",
    "00001000",
    "00000000",

-- 0x1e:
-- u+2339:
    "01111100",
    "01010100",
    "01000100",
    "01111100",
    "01000100",
    "01010100",
    "01111100",
    "00000000",

-- 0x1f:
-- u+2336:
    "00000000",
    "00000000",
    "01111100",
    "00010000",
    "00010000",
    "00010000",
    "01111100",
    "00000000",

-- # [ ] SPACE
-- 0x20:
-- u+0020:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",


-- # [!] EXCLAMATION MARK
-- 0x21:
-- u+0021:
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00000000",
    "00000000",
    "00001000",
    "00000000",


-- # ["] QUOTATION MARK
-- 0x22:
-- u+0022:
    "00100100",
    "00100100",
    "00100100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",


-- # [-- #] NUMBER SIGN
-- 0x23:
-- u+0023:
    "00100100",
    "00100100",
    "01111110",
    "00100100",
    "01111110",
    "00100100",
    "00100100",
    "00000000",


-- # [$] DOLLAR SIGN
-- 0x24:
-- u+0024:
    "00001000",
    "00011110",
    "00101000",
    "00011100",
    "00001010",
    "00111100",
    "00001000",
    "00000000",


-- # [%] PERCENT SIGN
-- 0x25:
-- u+0025:
    "00000000",
    "01100010",
    "01100100",
    "00001000",
    "00010000",
    "00100110",
    "01000110",
    "00000000",


-- # [&] AMPERSAND
-- 0x26:
-- u+0026:
    "00110000",
    "01001000",
    "01001000",
    "00110000",
    "01001010",
    "01000100",
    "00111010",
    "00000000",


-- # ['] APOSTROPHE
-- 0x27:
-- u+0027:
    "00000100",
    "00001000",
    "00010000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",


-- # [(] LEFT PARENTHESIS
-- 0x28:
-- u+0028:
    "00000100",
    "00001000",
    "00010000",
    "00010000",
    "00010000",
    "00001000",
    "00000100",
    "00000000",


-- # [)] RIGHT PARENTHESIS
-- 0x29:
-- u+0029:
    "00100000",
    "00010000",
    "00001000",
    "00001000",
    "00001000",
    "00010000",
    "00100000",
    "00000000",


-- # [*] ASTERISK
-- 0x2a:
-- u+002a:
    "00001000",
    "00101010",
    "00011100",
    "00111110",
    "00011100",
    "00101010",
    "00001000",
    "00000000",


-- # [+] PLUS SIGN
-- 0x2b:
-- u+002b:
    "00000000",
    "00001000",
    "00001000",
    "00111110",
    "00001000",
    "00001000",
    "00000000",
    "00000000",


-- # [,] COMMA
-- 0x2c:
-- u+002c:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00001000",
    "00001000",
    "00010000",


-- # [-] HYPHEN-MINUS
-- 0x2d:
-- u+002d:
    "00000000",
    "00000000",
    "00000000",
    "01111110",
    "00000000",
    "00000000",
    "00000000",
    "00000000",


-- # [0] FULL STOP
-- 0x2e:
-- u+002e:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00011000",
    "00011000",
    "00000000",


-- # [/] SOLIDUS
-- 0x2f:
-- u+002f:
    "00000000",
    "00000010",
    "00000100",
    "00001000",
    "00010000",
    "00100000",
    "01000000",
    "00000000",


-- # [0] DIGIT ZERO
-- 0x30:
-- u+0030:
    "00111100",
    "01000010",
    "01000110",
    "01011010",
    "01100010",
    "01000010",
    "00111100",
    "00000000",


-- # [1] DIGIT ONE
-- 0x31:
-- u+0031:
    "00001000",
    "00011000",
    "00101000",
    "00001000",
    "00001000",
    "00001000",
    "00111110",
    "00000000",


-- # [2] DIGIT TWO
-- 0x32:
-- u+0032:
    "00111100",
    "01000010",
    "00000010",
    "00001100",
    "00110000",
    "01000000",
    "01111110",
    "00000000",


-- # [3] DIGIT THREE
-- 0x33:
-- u+0033:
    "00111100",
    "01000010",
    "00000010",
    "00011100",
    "00000010",
    "01000010",
    "00111100",
    "00000000",


-- # [4] DIGIT FOUR
-- 0x34:
-- u+0034:
    "00000100",
    "00001100",
    "00010100",
    "00100100",
    "01111110",
    "00000100",
    "00000100",
    "00000000",


-- # [5] DIGIT FIVE
-- 0x35:
-- u+0035:
    "01111110",
    "01000000",
    "01111000",
    "00000100",
    "00000010",
    "01000100",
    "00111000",
    "00000000",


-- # [6] DIGIT SIX
-- 0x36:
-- u+0036:
    "00011100",
    "00100000",
    "01000000",
    "01111100",
    "01000010",
    "01000010",
    "00111100",
    "00000000",


-- # [7] DIGIT SEVEN
-- 0x37:
-- u+0037:
    "01111110",
    "01000010",
    "00000100",
    "00001000",
    "00010000",
    "00010000",
    "00010000",
    "00000000",


-- # [8] DIGIT EIGHT
-- 0x38:
-- u+0038:
    "00111100",
    "01000010",
    "01000010",
    "00111100",
    "01000010",
    "01000010",
    "00111100",
    "00000000",


-- # [9] DIGIT NINE
-- 0x39:
-- u+0039:
    "00111100",
    "01000010",
    "01000010",
    "00111110",
    "00000010",
    "00000100",
    "00111000",
    "00000000",


-- # [:] COLON
-- 0x3a:
-- u+003a:
    "00000000",
    "00000000",
    "00001000",
    "00000000",
    "00000000",
    "00001000",
    "00000000",
    "00000000",


-- # [;] SEMICOLON
-- 0x3b:
-- u+003b:
    "00000000",
    "00000000",
    "00001000",
    "00000000",
    "00000000",
    "00001000",
    "00001000",
    "00010000",


-- # [<] LESS-THAN SIGN
-- 0x3c:
-- u+003c:
    "00001110",
    "00011000",
    "00110000",
    "01100000",
    "00110000",
    "00011000",
    "00001110",
    "00000000",


-- # [=] EQUALS SIGN
-- 0x3d:
-- u+003d:
    "00000000",
    "00000000",
    "01111110",
    "00000000",
    "01111110",
    "00000000",
    "00000000",
    "00000000",


-- # [>] GREATER-THAN SIGN
-- 0x3e:
-- u+003e:
    "01110000",
    "00011000",
    "00001100",
    "00000110",
    "00001100",
    "00011000",
    "01110000",
    "00000000",


-- # [?] QUESTION MARK
-- 0x3f:
-- u+003f:
    "00111100",
    "01000010",
    "00000010",
    "00001100",
    "00010000",
    "00000000",
    "00010000",
    "00000000",


-- # [1] COMMERCIAL AT
-- 0x40:
-- u+0040:
    "00011100",
    "00100010",
    "01001010",
    "01010110",
    "01001100",
    "00100000",
    "00011110",
    "00000000",


-- # [A] LATIN CAPITAL LETTER A
-- 0x41:
-- u+0041:
    "00011000",
    "00100100",
    "01000010",
    "01111110",
    "01000010",
    "01000010",
    "01000010",
    "00000000",


-- # [B] LATIN CAPITAL LETTER B
-- 0x42:
-- u+0042:
    "01111100",
    "00100010",
    "00100010",
    "00111100",
    "00100010",
    "00100010",
    "01111100",
    "00000000",


-- # [C] LATIN CAPITAL LETTER C
-- 0x43:
-- u+0043:
    "00011100",
    "00100010",
    "01000000",
    "01000000",
    "01000000",
    "00100010",
    "00011100",
    "00000000",


-- # [D] LATIN CAPITAL LETTER D
-- 0x44:
-- u+0044:
    "01111000",
    "00100100",
    "00100010",
    "00100010",
    "00100010",
    "00100100",
    "01111000",
    "00000000",


-- # [E] LATIN CAPITAL LETTER E
-- 0x45:
-- u+0045:
    "01111110",
    "01000000",
    "01000000",
    "01111000",
    "01000000",
    "01000000",
    "01111110",
    "00000000",


-- # [F] LATIN CAPITAL LETTER F
-- 0x46:
-- u+0046:
    "01111110",
    "01000000",
    "01000000",
    "01111000",
    "01000000",
    "01000000",
    "01000000",
    "00000000",


-- # [G] LATIN CAPITAL LETTER G
-- 0x47:
-- u+0047:
    "00011100",
    "00100010",
    "01000000",
    "01001110",
    "01000010",
    "00100010",
    "00011100",
    "00000000",


-- # [H] LATIN CAPITAL LETTER H
-- 0x48:
-- u+0048:
    "01000010",
    "01000010",
    "01000010",
    "01111110",
    "01000010",
    "01000010",
    "01000010",
    "00000000",


-- # [I] LATIN CAPITAL LETTER I
-- 0x49:
-- u+0049:
    "00011100",
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00011100",
    "00000000",


-- # [J] LATIN CAPITAL LETTER J
-- 0x4a:
-- u+004a:
    "00001110",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "01000100",
    "00111000",
    "00000000",


-- # [K] LATIN CAPITAL LETTER K
-- 0x4b:
-- u+004b:
    "01000010",
    "01000100",
    "01001000",
    "01110000",
    "01001000",
    "01000100",
    "01000010",
    "00000000",


-- # [L] LATIN CAPITAL LETTER L
-- 0x4c:
-- u+004c:
    "01000000",
    "01000000",
    "01000000",
    "01000000",
    "01000000",
    "01000000",
    "01111110",
    "00000000",


-- # [M] LATIN CAPITAL LETTER M
-- 0x4d:
-- u+004d:
    "01000010",
    "01100110",
    "01011010",
    "01011010",
    "01000010",
    "01000010",
    "01000010",
    "00000000",


-- # [N] LATIN CAPITAL LETTER N
-- 0x4e:
-- u+004e:
    "01000010",
    "01100010",
    "01010010",
    "01001010",
    "01000110",
    "01000010",
    "01000010",
    "00000000",


-- # [O] LATIN CAPITAL LETTER O
-- 0x4f:
-- u+004f:
    "00011000",
    "00100100",
    "01000010",
    "01000010",
    "01000010",
    "00100100",
    "00011000",
    "00000000",


-- # [P] LATIN CAPITAL LETTER P
-- 0x50:
-- u+0050:
    "01111100",
    "01000010",
    "01000010",
    "01111100",
    "01000000",
    "01000000",
    "01000000",
    "00000000",


-- # [Q] LATIN CAPITAL LETTER Q
-- 0x51:
-- u+0051:
    "00011000",
    "00100100",
    "01000010",
    "01000010",
    "01001010",
    "00100100",
    "00011010",
    "00000000",


-- # [R] LATIN CAPITAL LETTER R
-- 0x52:
-- u+0052:
    "01111100",
    "01000010",
    "01000010",
    "01111100",
    "01001000",
    "01000100",
    "01000010",
    "00000000",


-- # [S] LATIN CAPITAL LETTER S
-- 0x53:
-- u+0053:
    "00111100",
    "01000010",
    "01000000",
    "00111100",
    "00000010",
    "01000010",
    "00111100",
    "00000000",


-- # [T] LATIN CAPITAL LETTER T
-- 0x54:
-- u+0054:
    "00111110",
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00000000",


-- # [U] LATIN CAPITAL LETTER U
-- 0x55:
-- u+0055:
    "01000010",
    "01000010",
    "01000010",
    "01000010",
    "01000010",
    "01000010",
    "00111100",
    "00000000",


-- # [V] LATIN CAPITAL LETTER V
-- 0x56:
-- u+0056:
    "01000010",
    "01000010",
    "01000010",
    "00100100",
    "00100100",
    "00011000",
    "00011000",
    "00000000",


-- # [W] LATIN CAPITAL LETTER W
-- 0x57:
-- u+0057:
    "01000010",
    "01000010",
    "01000010",
    "01011010",
    "01011010",
    "01100110",
    "01000010",
    "00000000",


-- # [X] LATIN CAPITAL LETTER X
-- 0x58:
-- u+0058:
    "01000010",
    "01000010",
    "00100100",
    "00011000",
    "00100100",
    "01000010",
    "01000010",
    "00000000",


-- # [Y] LATIN CAPITAL LETTER Y
-- 0x59:
-- u+0059:
    "00100010",
    "00100010",
    "00100010",
    "00011100",
    "00001000",
    "00001000",
    "00001000",
    "00000000",


-- # [Z] LATIN CAPITAL LETTER Z
-- 0x5a:
-- u+005a:
    "01111110",
    "00000010",
    "00000100",
    "00011000",
    "00100000",
    "01000000",
    "01111110",
    "00000000",


-- # [[] LEFT SQUARE BRACKET
-- 0x5b:
-- u+005b:
    "00111100",
    "00100000",
    "00100000",
    "00100000",
    "00100000",
    "00100000",
    "00111100",
    "00000000",


-- # [\] REVERSE SOLIDUS
-- 0x5c:
-- u+005c:
    "00000000",
    "01000000",
    "00100000",
    "00010000",
    "00001000",
    "00000100",
    "00000010",
    "00000000",


-- # []] RIGHT SQUARE BRACKET
-- 0x5d:
-- u+005d:
    "00111100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00000100",
    "00111100",
    "00000000",


-- # [^] CIRCUMFLEX ACCENT
-- 0x5e:
-- u+005e:
    "00010000",
    "00101000",
    "01000100",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",


-- # [_] LOW LINE
-- 0x5f:
-- u+005f:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "11111110",


-- # [`] GRAVE ACCENT
-- 0x60:
-- u+0060:
    "00100000",
    "00010000",
    "00001000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00000000",


-- # [a] LATIN SMALL LETTER A
-- 0x61:
-- u+0061:
    "00000000",
    "00000000",
    "00111000",
    "00000100",
    "00111100",
    "01000100",
    "00111010",
    "00000000",


-- # [b] LATIN SMALL LETTER B
-- 0x62:
-- u+0062:
    "01000000",
    "01000000",
    "01011100",
    "01100010",
    "01000010",
    "01100010",
    "01011100",
    "00000000",


-- # [c] LATIN SMALL LETTER C
-- 0x63:
-- u+0063:
    "00000000",
    "00000000",
    "00111100",
    "01000010",
    "01000000",
    "01000010",
    "00111100",
    "00000000",


-- # [d] LATIN SMALL LETTER D
-- 0x64:
-- u+0064:
    "00000010",
    "00000010",
    "00111010",
    "01000110",
    "01000010",
    "01000110",
    "00111010",
    "00000000",


-- # [e] LATIN SMALL LETTER E
-- 0x65:
-- u+0065:
    "00000000",
    "00000000",
    "00111100",
    "01000010",
    "01111110",
    "01000000",
    "00111100",
    "00000000",


-- # [f] LATIN SMALL LETTER F
-- 0x66:
-- u+0066:
    "00001100",
    "00010010",
    "00010000",
    "01111100",
    "00010000",
    "00010000",
    "00010000",
    "00000000",


-- # [g] LATIN SMALL LETTER G
-- 0x67:
-- u+0067:
    "00000000",
    "00000000",
    "00111010",
    "01000110",
    "01000110",
    "00111010",
    "00000010",
    "00111100",


-- # [h] LATIN SMALL LETTER H
-- 0x68:
-- u+0068:
    "01000000",
    "01000000",
    "01011100",
    "01100010",
    "01000010",
    "01000010",
    "01000010",
    "00000000",


-- # [i] LATIN SMALL LETTER I
-- 0x69:
-- u+0069:
    "00001000",
    "00000000",
    "00011000",
    "00001000",
    "00001000",
    "00001000",
    "00011100",
    "00000000",


-- # [j] LATIN SMALL LETTER J
-- 0x6a:
-- u+006a:
    "00000100",
    "00000000",
    "00001100",
    "00000100",
    "00000100",
    "00000100",
    "01000100",
    "00111000",


-- # [k] LATIN SMALL LETTER K
-- 0x6b:
-- u+006b:
    "01000000",
    "01000000",
    "01000100",
    "01001000",
    "01010000",
    "01101000",
    "01000100",
    "00000000",


-- # [l] LATIN SMALL LETTER L
-- 0x6c:
-- u+006c:
    "00011000",
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00011100",
    "00000000",


-- # [m] LATIN SMALL LETTER M
-- 0x6d:
-- u+006d:
    "00000000",
    "00000000",
    "01110110",
    "01001001",
    "01001001",
    "01001001",
    "01001001",
    "00000000",


-- # [n] LATIN SMALL LETTER N
-- 0x6e:
-- u+006e:
    "00000000",
    "00000000",
    "01011100",
    "01100010",
    "01000010",
    "01000010",
    "01000010",
    "00000000",


-- # [o] LATIN SMALL LETTER O
-- 0x6f:
-- u+006f:
    "00000000",
    "00000000",
    "00111100",
    "01000010",
    "01000010",
    "01000010",
    "00111100",
    "00000000",


-- # [p] LATIN SMALL LETTER P
-- 0x70:
-- u+0070:
    "00000000",
    "00000000",
    "01011100",
    "01100010",
    "01100010",
    "01011100",
    "01000000",
    "01000000",


-- # [q] LATIN SMALL LETTER Q
-- 0x71:
-- u+0071:
    "00000000",
    "00000000",
    "00111010",
    "01000110",
    "01000110",
    "00111010",
    "00000010",
    "00000010",


-- # [r] LATIN SMALL LETTER R
-- 0x72:
-- u+0072:
    "00000000",
    "00000000",
    "01011100",
    "01100010",
    "01000000",
    "01000000",
    "01000000",
    "00000000",


-- # [s] LATIN SMALL LETTER S
-- 0x73:
-- u+0073:
    "00000000",
    "00000000",
    "00111110",
    "01000000",
    "00111100",
    "00000010",
    "01111100",
    "00000000",


-- # [t] LATIN SMALL LETTER T
-- 0x74:
-- u+0074:
    "00010000",
    "00010000",
    "01111100",
    "00010000",
    "00010000",
    "00010010",
    "00001100",
    "00000000",


-- # [u] LATIN SMALL LETTER U
-- 0x75:
-- u+0075:
    "00000000",
    "00000000",
    "01000010",
    "01000010",
    "01000010",
    "01000110",
    "00111010",
    "00000000",


-- # [v] LATIN SMALL LETTER V
-- 0x76:
-- u+0076:
    "00000000",
    "00000000",
    "01000010",
    "01000010",
    "01000010",
    "00100100",
    "00011000",
    "00000000",


-- # [w] LATIN SMALL LETTER W
-- 0x77:
-- u+0077:
    "00000000",
    "00000000",
    "01000001",
    "01001001",
    "01001001",
    "01001001",
    "00110110",
    "00000000",


-- # [x] LATIN SMALL LETTER X
-- 0x78:
-- u+0078:
    "00000000",
    "00000000",
    "01000010",
    "00100100",
    "00011000",
    "00100100",
    "01000010",
    "00000000",


-- # [y] LATIN SMALL LETTER Y
-- 0x79:
-- u+0079:
    "00000000",
    "00000000",
    "01000010",
    "01000010",
    "01000110",
    "00111010",
    "00000010",
    "00111100",


-- # [z] LATIN SMALL LETTER Z
-- 0x7a:
-- u+007a:
    "00000000",
    "00000000",
    "01111110",
    "00000100",
    "00011000",
    "00100000",
    "01111110",
    "00000000",


-- # [{] LEFT CURLY BRACKET
-- 0x7b:
-- u+007b:
    "00011000",
    "00100000",
    "00100000",
    "01000000",
    "00100000",
    "00100000",
    "00011000",
    "00000000",


-- # [|] VERTICAL LINE
-- 0x7c:
-- u+007c:
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00001000",
    "00001000",


-- # [}] RIGHT CURLY BRACKET
-- 0x7d:
-- u+007d:
    "00110000",
    "00001000",
    "00001000",
    "00000100",
    "00001000",
    "00001000",
    "00110000",
    "00000000",


-- # [~] TILDE
-- 0x7e:
-- u+007e:
    "00000000",
    "00000000",
    "00000000",
    "00100000",
    "01010100",
    "00001000",
    "00000000",
    "00000000",

-- 0x7f:
    "00000000",
    "00000000",
    "00000000",
    "00000000",
    "00111110",
    "00111110",
    "00111110",
    "00111110"
    );
begin

    dataOut <= ROM(to_integer(unsigned(addrIn)));

end architecture rtl;